MACRO tt_um_jnw_wulffern
  CLASS BLOCK ;
  FOREIGN tt_um_jnw_wulffern ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 10.020 204.890 17.620 210.170 ;
        RECT 19.020 204.390 26.620 209.670 ;
        RECT 28.020 204.390 35.620 209.670 ;
        RECT 37.020 204.390 44.620 209.670 ;
        RECT 55.020 204.390 62.620 209.670 ;
        RECT 73.420 204.390 81.020 209.670 ;
        RECT 82.420 204.390 90.020 209.670 ;
        RECT 91.420 204.390 99.020 209.670 ;
        RECT 100.420 204.890 108.020 210.170 ;
        RECT 10.020 197.390 17.620 202.670 ;
        RECT 19.020 197.390 26.620 202.670 ;
        RECT 28.020 197.390 35.620 202.670 ;
        RECT 37.020 197.390 44.620 202.670 ;
        RECT 46.020 197.390 53.620 202.670 ;
        RECT 55.020 197.390 62.620 202.670 ;
        RECT 64.420 197.390 72.020 202.670 ;
        RECT 73.420 197.390 81.020 202.670 ;
        RECT 82.420 197.390 90.020 202.670 ;
        RECT 91.420 197.390 99.020 202.670 ;
        RECT 100.420 197.390 108.020 202.670 ;
      LAYER pwell ;
        RECT 110.840 195.790 116.600 210.190 ;
      LAYER nwell ;
        RECT 10.020 190.390 17.620 195.670 ;
        RECT 19.020 190.390 26.620 195.670 ;
        RECT 28.020 190.390 35.620 195.670 ;
        RECT 37.020 190.390 44.620 195.670 ;
        RECT 55.020 190.390 62.620 195.670 ;
        RECT 73.420 190.390 81.020 195.670 ;
        RECT 82.420 190.390 90.020 195.670 ;
        RECT 91.420 190.390 99.020 195.670 ;
        RECT 100.420 190.390 108.020 195.670 ;
      LAYER pwell ;
        RECT 14.840 172.790 33.560 187.190 ;
      LAYER nwell ;
        RECT 37.020 181.890 44.620 187.170 ;
        RECT 46.020 181.390 53.620 186.670 ;
        RECT 64.420 181.390 72.020 186.670 ;
        RECT 73.420 181.890 81.020 187.170 ;
        RECT 37.020 174.390 44.620 179.670 ;
        RECT 46.020 174.390 53.620 179.670 ;
        RECT 64.420 174.390 72.020 179.670 ;
        RECT 73.420 174.390 81.020 179.670 ;
      LAYER pwell ;
        RECT 84.480 172.790 103.200 187.190 ;
        RECT 110.840 177.790 116.600 192.190 ;
        RECT 14.840 154.790 33.560 169.190 ;
        RECT 37.020 161.390 44.620 171.670 ;
        RECT 46.020 161.390 53.620 171.670 ;
        RECT 64.420 161.390 72.020 171.670 ;
        RECT 73.420 161.390 81.020 171.670 ;
        RECT 38.020 157.325 44.720 158.090 ;
        RECT 38.020 152.155 38.785 157.325 ;
        RECT 43.955 152.155 44.720 157.325 ;
        RECT 38.020 151.390 44.720 152.155 ;
        RECT 46.020 157.325 52.720 158.090 ;
        RECT 46.020 152.155 46.785 157.325 ;
        RECT 51.955 152.155 52.720 157.325 ;
        RECT 46.020 151.390 52.720 152.155 ;
        RECT 54.020 157.325 60.720 158.090 ;
        RECT 54.020 152.155 54.785 157.325 ;
        RECT 59.955 152.155 60.720 157.325 ;
      LAYER nwell ;
        RECT 62.820 155.790 68.520 159.390 ;
      LAYER pwell ;
        RECT 68.520 155.790 74.220 159.390 ;
        RECT 84.480 154.790 103.200 169.190 ;
        RECT 110.840 159.790 116.600 174.190 ;
        RECT 54.020 151.390 60.720 152.155 ;
        RECT 14.840 136.790 33.560 151.190 ;
        RECT 38.020 149.325 44.720 150.090 ;
        RECT 38.020 144.155 38.785 149.325 ;
        RECT 43.955 144.155 44.720 149.325 ;
        RECT 38.020 143.390 44.720 144.155 ;
        RECT 46.020 149.325 52.720 150.090 ;
        RECT 46.020 144.155 46.785 149.325 ;
        RECT 51.955 144.155 52.720 149.325 ;
        RECT 46.020 143.390 52.720 144.155 ;
        RECT 54.020 149.325 60.720 150.090 ;
        RECT 54.020 144.155 54.785 149.325 ;
        RECT 59.955 144.155 60.720 149.325 ;
        RECT 54.020 143.390 60.720 144.155 ;
        RECT 38.020 141.325 44.720 142.090 ;
        RECT 38.020 136.155 38.785 141.325 ;
        RECT 43.955 136.155 44.720 141.325 ;
        RECT 38.020 135.390 44.720 136.155 ;
        RECT 46.020 141.325 52.720 142.090 ;
        RECT 46.020 136.155 46.785 141.325 ;
        RECT 51.955 136.155 52.720 141.325 ;
        RECT 46.020 135.390 52.720 136.155 ;
        RECT 54.020 141.325 60.720 142.090 ;
        RECT 54.020 136.155 54.785 141.325 ;
        RECT 59.955 136.155 60.720 141.325 ;
        RECT 54.020 135.390 60.720 136.155 ;
        RECT 62.020 133.970 67.720 154.290 ;
        RECT 59.520 133.890 67.720 133.970 ;
      LAYER nwell ;
        RECT 67.720 133.890 73.420 154.290 ;
      LAYER pwell ;
        RECT 110.840 141.790 116.600 156.190 ;
        RECT 14.840 118.790 33.560 133.190 ;
        RECT 38.840 118.790 57.560 133.190 ;
        RECT 59.520 123.890 66.480 133.890 ;
      LAYER li1 ;
        RECT 10.520 210.870 107.520 211.890 ;
        RECT 109.020 210.950 119.020 211.890 ;
        RECT 10.460 209.910 107.580 210.870 ;
        RECT 10.460 190.870 11.420 209.910 ;
        RECT 12.380 208.930 14.620 209.330 ;
        RECT 11.740 206.930 12.060 208.130 ;
        RECT 13.020 207.330 15.260 207.730 ;
        RECT 15.580 206.930 15.900 208.130 ;
        RECT 12.380 205.730 14.620 206.130 ;
        RECT 12.380 201.430 14.620 201.830 ;
        RECT 11.740 199.430 12.060 200.630 ;
        RECT 13.020 199.830 15.260 200.230 ;
        RECT 15.580 199.430 15.900 200.630 ;
        RECT 12.380 198.230 14.620 198.630 ;
        RECT 12.380 194.430 14.620 194.830 ;
        RECT 11.740 192.430 12.060 193.630 ;
        RECT 13.020 192.830 15.260 193.230 ;
        RECT 15.580 192.430 15.900 193.630 ;
        RECT 12.380 191.230 14.620 191.630 ;
        RECT 16.220 190.870 20.420 209.910 ;
        RECT 21.380 208.430 23.620 208.830 ;
        RECT 20.740 206.430 21.060 207.630 ;
        RECT 22.020 206.830 24.260 207.230 ;
        RECT 24.580 206.430 24.900 207.630 ;
        RECT 21.380 205.230 23.620 205.630 ;
        RECT 21.380 201.430 23.620 201.830 ;
        RECT 20.740 199.430 21.060 200.630 ;
        RECT 22.020 199.830 24.260 200.230 ;
        RECT 24.580 199.430 24.900 200.630 ;
        RECT 21.380 198.230 23.620 198.630 ;
        RECT 21.380 194.430 23.620 194.830 ;
        RECT 20.740 192.430 21.060 193.630 ;
        RECT 22.020 192.830 24.260 193.230 ;
        RECT 24.580 192.430 24.900 193.630 ;
        RECT 21.380 191.230 23.620 191.630 ;
        RECT 25.220 190.870 29.420 209.910 ;
        RECT 30.380 208.430 32.620 208.830 ;
        RECT 29.740 206.430 30.060 207.630 ;
        RECT 31.020 206.830 33.260 207.230 ;
        RECT 33.580 206.430 33.900 207.630 ;
        RECT 30.380 205.230 32.620 205.630 ;
        RECT 30.380 201.430 32.620 201.830 ;
        RECT 29.740 199.430 30.060 200.630 ;
        RECT 31.020 199.830 33.260 200.230 ;
        RECT 33.580 199.430 33.900 200.630 ;
        RECT 30.380 198.230 32.620 198.630 ;
        RECT 30.380 194.430 32.620 194.830 ;
        RECT 29.740 192.430 30.060 193.630 ;
        RECT 31.020 192.830 33.260 193.230 ;
        RECT 33.580 192.430 33.900 193.630 ;
        RECT 30.380 191.230 32.620 191.630 ;
        RECT 34.220 190.870 38.420 209.910 ;
        RECT 39.380 208.430 41.620 208.830 ;
        RECT 38.740 206.430 39.060 207.630 ;
        RECT 40.020 206.830 42.260 207.230 ;
        RECT 42.580 206.430 42.900 207.630 ;
        RECT 39.380 205.230 41.620 205.630 ;
        RECT 43.220 202.410 56.420 209.910 ;
        RECT 57.380 208.430 59.620 208.830 ;
        RECT 56.740 206.430 57.060 207.630 ;
        RECT 58.020 206.830 60.260 207.230 ;
        RECT 60.580 206.430 60.900 207.630 ;
        RECT 57.380 205.230 59.620 205.630 ;
        RECT 39.380 201.430 41.620 201.830 ;
        RECT 38.740 199.430 39.060 200.630 ;
        RECT 40.020 199.830 42.260 200.230 ;
        RECT 42.580 199.430 42.900 200.630 ;
        RECT 39.380 198.230 41.620 198.630 ;
        RECT 43.220 197.870 47.420 202.410 ;
        RECT 48.380 201.430 50.620 201.830 ;
        RECT 47.740 199.430 48.060 200.630 ;
        RECT 49.020 199.830 51.260 200.230 ;
        RECT 51.580 199.430 51.900 200.630 ;
        RECT 48.380 198.230 50.620 198.630 ;
        RECT 52.220 197.870 56.420 202.410 ;
        RECT 61.220 202.410 74.820 209.910 ;
        RECT 76.420 208.430 78.660 208.830 ;
        RECT 75.140 206.430 75.460 207.630 ;
        RECT 75.780 206.830 78.020 207.230 ;
        RECT 78.980 206.430 79.300 207.630 ;
        RECT 76.420 205.230 78.660 205.630 ;
        RECT 57.380 201.430 59.620 201.830 ;
        RECT 56.740 199.430 57.060 200.630 ;
        RECT 58.020 199.830 60.260 200.230 ;
        RECT 60.580 199.430 60.900 200.630 ;
        RECT 57.380 198.230 59.620 198.630 ;
        RECT 39.380 194.430 41.620 194.830 ;
        RECT 38.740 192.430 39.060 193.630 ;
        RECT 40.020 192.830 42.260 193.230 ;
        RECT 42.580 192.430 42.900 193.630 ;
        RECT 39.380 191.230 41.620 191.630 ;
        RECT 43.220 190.870 56.420 197.870 ;
        RECT 61.220 197.870 65.820 202.410 ;
        RECT 67.420 201.430 69.660 201.830 ;
        RECT 66.140 199.430 66.460 200.630 ;
        RECT 66.780 199.830 69.020 200.230 ;
        RECT 69.980 199.430 70.300 200.630 ;
        RECT 67.420 198.230 69.660 198.630 ;
        RECT 70.620 197.870 74.820 202.410 ;
        RECT 76.420 201.430 78.660 201.830 ;
        RECT 75.140 199.430 75.460 200.630 ;
        RECT 75.780 199.830 78.020 200.230 ;
        RECT 78.980 199.430 79.300 200.630 ;
        RECT 76.420 198.230 78.660 198.630 ;
        RECT 57.380 194.430 59.620 194.830 ;
        RECT 56.740 192.430 57.060 193.630 ;
        RECT 58.020 192.830 60.260 193.230 ;
        RECT 60.580 192.430 60.900 193.630 ;
        RECT 57.380 191.230 59.620 191.630 ;
        RECT 61.220 190.870 74.820 197.870 ;
        RECT 76.420 194.430 78.660 194.830 ;
        RECT 75.140 192.430 75.460 193.630 ;
        RECT 75.780 192.830 78.020 193.230 ;
        RECT 78.980 192.430 79.300 193.630 ;
        RECT 76.420 191.230 78.660 191.630 ;
        RECT 79.620 190.870 83.820 209.910 ;
        RECT 85.420 208.430 87.660 208.830 ;
        RECT 84.140 206.430 84.460 207.630 ;
        RECT 84.780 206.830 87.020 207.230 ;
        RECT 87.980 206.430 88.300 207.630 ;
        RECT 85.420 205.230 87.660 205.630 ;
        RECT 85.420 201.430 87.660 201.830 ;
        RECT 84.140 199.430 84.460 200.630 ;
        RECT 84.780 199.830 87.020 200.230 ;
        RECT 87.980 199.430 88.300 200.630 ;
        RECT 85.420 198.230 87.660 198.630 ;
        RECT 85.420 194.430 87.660 194.830 ;
        RECT 84.140 192.430 84.460 193.630 ;
        RECT 84.780 192.830 87.020 193.230 ;
        RECT 87.980 192.430 88.300 193.630 ;
        RECT 85.420 191.230 87.660 191.630 ;
        RECT 88.620 190.870 92.820 209.910 ;
        RECT 94.420 208.430 96.660 208.830 ;
        RECT 93.140 206.430 93.460 207.630 ;
        RECT 93.780 206.830 96.020 207.230 ;
        RECT 96.980 206.430 97.300 207.630 ;
        RECT 94.420 205.230 96.660 205.630 ;
        RECT 94.420 201.430 96.660 201.830 ;
        RECT 93.140 199.430 93.460 200.630 ;
        RECT 93.780 199.830 96.020 200.230 ;
        RECT 96.980 199.430 97.300 200.630 ;
        RECT 94.420 198.230 96.660 198.630 ;
        RECT 94.420 194.430 96.660 194.830 ;
        RECT 93.140 192.430 93.460 193.630 ;
        RECT 93.780 192.830 96.020 193.230 ;
        RECT 96.980 192.430 97.300 193.630 ;
        RECT 94.420 191.230 96.660 191.630 ;
        RECT 97.620 190.870 101.820 209.910 ;
        RECT 103.420 208.930 105.660 209.330 ;
        RECT 102.140 206.930 102.460 208.130 ;
        RECT 102.780 207.330 105.020 207.730 ;
        RECT 105.980 206.930 106.300 208.130 ;
        RECT 103.420 205.730 105.660 206.130 ;
        RECT 103.420 201.430 105.660 201.830 ;
        RECT 102.140 199.430 102.460 200.630 ;
        RECT 102.780 199.830 105.020 200.230 ;
        RECT 105.980 199.430 106.300 200.630 ;
        RECT 103.420 198.230 105.660 198.630 ;
        RECT 103.420 194.430 105.660 194.830 ;
        RECT 102.140 192.430 102.460 193.630 ;
        RECT 102.780 192.830 105.020 193.230 ;
        RECT 105.980 192.430 106.300 193.630 ;
        RECT 103.420 191.230 105.660 191.630 ;
        RECT 106.620 190.870 107.580 209.910 ;
        RECT 10.460 189.910 107.580 190.870 ;
        RECT 109.020 195.030 109.660 210.950 ;
        RECT 110.840 208.990 112.280 210.190 ;
        RECT 111.920 205.390 112.280 208.990 ;
        RECT 113.000 208.990 114.440 210.190 ;
        RECT 113.000 205.390 113.360 208.990 ;
        RECT 114.080 205.390 114.440 208.990 ;
        RECT 115.160 208.990 116.600 210.190 ;
        RECT 115.160 205.390 115.520 208.990 ;
        RECT 111.920 195.790 113.360 198.190 ;
        RECT 114.080 195.790 115.520 198.190 ;
        RECT 117.780 195.030 119.020 210.950 ;
        RECT 109.020 192.950 119.020 195.030 ;
        RECT 43.520 189.890 56.020 189.910 ;
        RECT 61.520 189.890 74.020 189.910 ;
        RECT 13.020 187.890 35.520 188.890 ;
        RECT 13.020 172.030 13.660 187.890 ;
        RECT 14.840 185.990 16.280 187.190 ;
        RECT 15.920 182.390 16.280 185.990 ;
        RECT 17.000 185.990 18.440 187.190 ;
        RECT 17.000 182.390 17.360 185.990 ;
        RECT 18.080 182.390 18.440 185.990 ;
        RECT 19.160 185.990 20.600 187.190 ;
        RECT 19.160 182.390 19.520 185.990 ;
        RECT 20.240 182.390 20.600 185.990 ;
        RECT 21.320 185.990 22.760 187.190 ;
        RECT 21.320 182.390 21.680 185.990 ;
        RECT 22.400 182.390 22.760 185.990 ;
        RECT 23.480 185.990 24.920 187.190 ;
        RECT 23.480 182.390 23.840 185.990 ;
        RECT 24.560 182.390 24.920 185.990 ;
        RECT 25.640 185.990 27.080 187.190 ;
        RECT 25.640 182.390 26.000 185.990 ;
        RECT 26.720 182.390 27.080 185.990 ;
        RECT 27.800 185.990 29.240 187.190 ;
        RECT 27.800 182.390 28.160 185.990 ;
        RECT 28.880 182.390 29.240 185.990 ;
        RECT 29.960 185.990 31.400 187.190 ;
        RECT 29.960 182.390 30.320 185.990 ;
        RECT 31.040 182.390 31.400 185.990 ;
        RECT 32.120 185.990 33.560 187.190 ;
        RECT 32.120 182.390 32.480 185.990 ;
        RECT 15.920 172.790 17.360 175.190 ;
        RECT 18.080 172.790 19.520 175.190 ;
        RECT 20.240 172.790 21.680 175.190 ;
        RECT 22.400 172.790 23.840 175.190 ;
        RECT 24.560 172.790 26.000 175.190 ;
        RECT 26.720 172.790 28.160 175.190 ;
        RECT 28.880 172.790 30.320 175.190 ;
        RECT 31.040 172.790 32.480 175.190 ;
        RECT 34.740 172.870 35.520 187.890 ;
        RECT 82.740 188.390 104.940 188.510 ;
        RECT 109.020 188.390 109.660 192.950 ;
        RECT 110.840 190.990 112.280 192.190 ;
        RECT 82.740 187.950 109.660 188.390 ;
        RECT 37.460 186.910 53.180 187.870 ;
        RECT 37.460 174.870 38.420 186.910 ;
        RECT 39.380 185.930 41.620 186.330 ;
        RECT 38.740 183.930 39.060 185.130 ;
        RECT 40.020 184.330 42.260 184.730 ;
        RECT 42.580 183.930 42.900 185.130 ;
        RECT 39.380 182.730 41.620 183.130 ;
        RECT 39.380 178.430 41.620 178.830 ;
        RECT 38.740 176.430 39.060 177.630 ;
        RECT 40.020 176.830 42.260 177.230 ;
        RECT 42.580 176.430 42.900 177.630 ;
        RECT 39.380 175.230 41.620 175.630 ;
        RECT 43.220 174.870 47.420 186.910 ;
        RECT 48.380 185.430 50.620 185.830 ;
        RECT 47.740 183.430 48.060 184.630 ;
        RECT 49.020 183.830 51.260 184.230 ;
        RECT 51.580 183.430 51.900 184.630 ;
        RECT 48.380 182.230 50.620 182.630 ;
        RECT 48.380 178.430 50.620 178.830 ;
        RECT 47.740 176.430 48.060 177.630 ;
        RECT 49.020 176.830 51.260 177.230 ;
        RECT 51.580 176.430 51.900 177.630 ;
        RECT 48.380 175.230 50.620 175.630 ;
        RECT 52.220 174.870 53.180 186.910 ;
        RECT 37.460 173.910 53.180 174.870 ;
        RECT 64.860 186.910 80.580 187.870 ;
        RECT 64.860 174.870 65.820 186.910 ;
        RECT 67.420 185.430 69.660 185.830 ;
        RECT 66.140 183.430 66.460 184.630 ;
        RECT 66.780 183.830 69.020 184.230 ;
        RECT 69.980 183.430 70.300 184.630 ;
        RECT 67.420 182.230 69.660 182.630 ;
        RECT 67.420 178.430 69.660 178.830 ;
        RECT 66.140 176.430 66.460 177.630 ;
        RECT 66.780 176.830 69.020 177.230 ;
        RECT 69.980 176.430 70.300 177.630 ;
        RECT 67.420 175.230 69.660 175.630 ;
        RECT 70.620 174.870 74.820 186.910 ;
        RECT 76.420 185.930 78.660 186.330 ;
        RECT 75.140 183.930 75.460 185.130 ;
        RECT 75.780 184.330 78.020 184.730 ;
        RECT 78.980 183.930 79.300 185.130 ;
        RECT 76.420 182.730 78.660 183.130 ;
        RECT 76.420 178.430 78.660 178.830 ;
        RECT 75.140 176.430 75.460 177.630 ;
        RECT 75.780 176.830 78.020 177.230 ;
        RECT 78.980 176.430 79.300 177.630 ;
        RECT 76.420 175.230 78.660 175.630 ;
        RECT 79.620 174.870 80.580 186.910 ;
        RECT 64.860 173.910 80.580 174.870 ;
        RECT 34.740 172.390 80.580 172.870 ;
        RECT 82.740 172.390 83.300 187.950 ;
        RECT 84.480 185.990 85.920 187.190 ;
        RECT 85.560 182.390 85.920 185.990 ;
        RECT 86.640 185.990 88.080 187.190 ;
        RECT 86.640 182.390 87.000 185.990 ;
        RECT 87.720 182.390 88.080 185.990 ;
        RECT 88.800 185.990 90.240 187.190 ;
        RECT 88.800 182.390 89.160 185.990 ;
        RECT 89.880 182.390 90.240 185.990 ;
        RECT 90.960 185.990 92.400 187.190 ;
        RECT 90.960 182.390 91.320 185.990 ;
        RECT 92.040 182.390 92.400 185.990 ;
        RECT 93.120 185.990 94.560 187.190 ;
        RECT 93.120 182.390 93.480 185.990 ;
        RECT 94.200 182.390 94.560 185.990 ;
        RECT 95.280 185.990 96.720 187.190 ;
        RECT 95.280 182.390 95.640 185.990 ;
        RECT 96.360 182.390 96.720 185.990 ;
        RECT 97.440 185.990 98.880 187.190 ;
        RECT 97.440 182.390 97.800 185.990 ;
        RECT 98.520 182.390 98.880 185.990 ;
        RECT 99.600 185.990 101.040 187.190 ;
        RECT 99.600 182.390 99.960 185.990 ;
        RECT 100.680 182.390 101.040 185.990 ;
        RECT 101.760 185.990 103.200 187.190 ;
        RECT 101.760 182.390 102.120 185.990 ;
        RECT 104.380 177.030 109.660 187.950 ;
        RECT 111.920 187.390 112.280 190.990 ;
        RECT 113.000 190.990 114.440 192.190 ;
        RECT 113.000 187.390 113.360 190.990 ;
        RECT 114.080 187.390 114.440 190.990 ;
        RECT 115.160 190.990 116.600 192.190 ;
        RECT 115.160 187.390 115.520 190.990 ;
        RECT 111.920 177.790 113.360 180.190 ;
        RECT 114.080 177.790 115.520 180.190 ;
        RECT 117.780 177.030 119.020 192.950 ;
        RECT 85.560 172.790 87.000 175.190 ;
        RECT 87.720 172.790 89.160 175.190 ;
        RECT 89.880 172.790 91.320 175.190 ;
        RECT 92.040 172.790 93.480 175.190 ;
        RECT 94.200 172.790 95.640 175.190 ;
        RECT 96.360 172.790 97.800 175.190 ;
        RECT 98.520 172.790 99.960 175.190 ;
        RECT 100.680 172.790 102.120 175.190 ;
        RECT 104.380 174.950 119.020 177.030 ;
        RECT 34.740 172.030 83.300 172.390 ;
        RECT 104.380 172.030 109.660 174.950 ;
        RECT 110.840 172.990 112.280 174.190 ;
        RECT 13.020 171.910 109.660 172.030 ;
        RECT 13.020 169.950 38.420 171.910 ;
        RECT 39.380 170.430 41.620 170.830 ;
        RECT 13.020 154.030 13.660 169.950 ;
        RECT 32.360 169.190 33.560 169.950 ;
        RECT 14.840 167.990 16.280 169.190 ;
        RECT 15.920 164.390 16.280 167.990 ;
        RECT 17.000 167.990 18.440 169.190 ;
        RECT 17.000 164.390 17.360 167.990 ;
        RECT 18.080 164.390 18.440 167.990 ;
        RECT 19.160 167.990 20.600 169.190 ;
        RECT 19.160 164.390 19.520 167.990 ;
        RECT 20.240 164.390 20.600 167.990 ;
        RECT 21.320 167.990 22.760 169.190 ;
        RECT 21.320 164.390 21.680 167.990 ;
        RECT 22.400 164.390 22.760 167.990 ;
        RECT 23.480 167.990 24.920 169.190 ;
        RECT 23.480 164.390 23.840 167.990 ;
        RECT 24.560 164.390 24.920 167.990 ;
        RECT 25.640 167.990 27.080 169.190 ;
        RECT 25.640 164.390 26.000 167.990 ;
        RECT 26.720 164.390 27.080 167.990 ;
        RECT 27.800 167.990 29.240 169.190 ;
        RECT 27.800 164.390 28.160 167.990 ;
        RECT 28.880 164.390 29.240 167.990 ;
        RECT 29.960 167.990 31.400 169.190 ;
        RECT 29.960 164.390 30.320 167.990 ;
        RECT 31.040 164.390 31.400 167.990 ;
        RECT 32.120 167.990 33.560 169.190 ;
        RECT 32.120 164.390 32.480 167.990 ;
        RECT 34.740 161.890 38.420 169.950 ;
        RECT 38.740 168.430 39.060 169.630 ;
        RECT 40.020 168.830 42.260 169.230 ;
        RECT 42.580 168.430 42.900 169.630 ;
        RECT 39.380 167.230 41.620 167.630 ;
        RECT 39.380 165.430 41.620 165.830 ;
        RECT 38.740 163.430 39.060 164.630 ;
        RECT 40.020 163.830 42.260 164.230 ;
        RECT 42.580 163.430 42.900 164.630 ;
        RECT 39.380 162.230 41.620 162.630 ;
        RECT 43.220 161.890 47.420 171.910 ;
        RECT 48.380 170.430 50.620 170.830 ;
        RECT 47.740 168.430 48.060 169.630 ;
        RECT 49.020 168.830 51.260 169.230 ;
        RECT 51.580 168.430 51.900 169.630 ;
        RECT 48.380 167.230 50.620 167.630 ;
        RECT 48.380 165.430 50.620 165.830 ;
        RECT 47.740 163.430 48.060 164.630 ;
        RECT 49.020 163.830 51.260 164.230 ;
        RECT 51.580 163.430 51.900 164.630 ;
        RECT 48.380 162.230 50.620 162.630 ;
        RECT 52.220 161.890 65.820 171.910 ;
        RECT 67.420 170.430 69.660 170.830 ;
        RECT 66.140 168.430 66.460 169.630 ;
        RECT 66.780 168.830 69.020 169.230 ;
        RECT 69.980 168.430 70.300 169.630 ;
        RECT 67.420 167.230 69.660 167.630 ;
        RECT 67.420 165.430 69.660 165.830 ;
        RECT 66.140 163.430 66.460 164.630 ;
        RECT 66.780 163.830 69.020 164.230 ;
        RECT 69.980 163.430 70.300 164.630 ;
        RECT 67.420 162.230 69.660 162.630 ;
        RECT 34.740 161.870 65.820 161.890 ;
        RECT 70.620 161.870 74.820 171.910 ;
        RECT 76.420 170.430 78.660 170.830 ;
        RECT 79.620 169.950 109.660 171.910 ;
        RECT 75.140 168.430 75.460 169.630 ;
        RECT 75.780 168.830 78.020 169.230 ;
        RECT 78.980 168.430 79.300 169.630 ;
        RECT 76.420 167.230 78.660 167.630 ;
        RECT 76.420 165.430 78.660 165.830 ;
        RECT 75.140 163.430 75.460 164.630 ;
        RECT 75.780 163.830 78.020 164.230 ;
        RECT 78.980 163.430 79.300 164.630 ;
        RECT 76.420 162.230 78.660 162.630 ;
        RECT 79.620 161.870 83.300 169.950 ;
        RECT 84.480 169.190 85.680 169.950 ;
        RECT 84.480 167.990 85.920 169.190 ;
        RECT 85.560 164.390 85.920 167.990 ;
        RECT 86.640 167.990 88.080 169.190 ;
        RECT 86.640 164.390 87.000 167.990 ;
        RECT 87.720 164.390 88.080 167.990 ;
        RECT 88.800 167.990 90.240 169.190 ;
        RECT 88.800 164.390 89.160 167.990 ;
        RECT 89.880 164.390 90.240 167.990 ;
        RECT 90.960 167.990 92.400 169.190 ;
        RECT 90.960 164.390 91.320 167.990 ;
        RECT 92.040 164.390 92.400 167.990 ;
        RECT 93.120 167.990 94.560 169.190 ;
        RECT 93.120 164.390 93.480 167.990 ;
        RECT 94.200 164.390 94.560 167.990 ;
        RECT 95.280 167.990 96.720 169.190 ;
        RECT 95.280 164.390 95.640 167.990 ;
        RECT 96.360 164.390 96.720 167.990 ;
        RECT 97.440 167.990 98.880 169.190 ;
        RECT 97.440 164.390 97.800 167.990 ;
        RECT 98.520 164.390 98.880 167.990 ;
        RECT 99.600 167.990 101.040 169.190 ;
        RECT 99.600 164.390 99.960 167.990 ;
        RECT 100.680 164.390 101.040 167.990 ;
        RECT 101.760 167.990 103.200 169.190 ;
        RECT 101.760 164.390 102.120 167.990 ;
        RECT 34.740 160.910 83.300 161.870 ;
        RECT 34.740 160.390 65.520 160.910 ;
        RECT 15.920 154.790 17.360 157.190 ;
        RECT 18.080 154.790 19.520 157.190 ;
        RECT 20.240 154.790 21.680 157.190 ;
        RECT 22.400 154.790 23.840 157.190 ;
        RECT 24.560 154.790 26.000 157.190 ;
        RECT 26.720 154.790 28.160 157.190 ;
        RECT 28.880 154.790 30.320 157.190 ;
        RECT 31.040 154.790 32.480 157.190 ;
        RECT 34.740 156.785 61.020 160.390 ;
        RECT 63.120 157.770 64.020 158.990 ;
        RECT 65.970 158.240 70.320 158.540 ;
        RECT 64.920 157.840 65.820 158.140 ;
        RECT 71.220 157.840 72.120 158.140 ;
        RECT 61.940 156.810 64.020 157.770 ;
        RECT 66.780 157.740 67.620 157.760 ;
        RECT 69.480 157.740 70.320 157.760 ;
        RECT 66.720 157.440 67.620 157.740 ;
        RECT 69.420 157.440 70.320 157.740 ;
        RECT 70.620 157.540 71.520 157.840 ;
        RECT 73.020 157.730 73.920 158.990 ;
        RECT 64.920 157.040 65.820 157.340 ;
        RECT 70.620 157.240 70.920 157.540 ;
        RECT 70.020 156.940 70.920 157.240 ;
        RECT 71.220 157.040 72.570 157.340 ;
        RECT 34.740 154.030 39.325 156.785 ;
        RECT 13.020 152.695 39.325 154.030 ;
        RECT 39.635 153.005 43.105 156.475 ;
        RECT 43.415 152.695 47.325 156.785 ;
        RECT 47.635 153.005 51.105 156.475 ;
        RECT 51.415 152.695 55.325 156.785 ;
        RECT 55.635 153.005 59.105 156.475 ;
        RECT 59.415 154.390 61.020 156.785 ;
        RECT 63.120 156.190 64.020 156.810 ;
        RECT 66.720 156.640 70.320 156.940 ;
        RECT 73.020 156.850 75.160 157.730 ;
        RECT 73.020 156.190 73.920 156.850 ;
        RECT 74.280 155.450 75.160 156.850 ;
        RECT 59.415 153.890 63.020 154.390 ;
        RECT 59.415 152.695 63.220 153.890 ;
        RECT 67.870 153.440 68.170 154.040 ;
        RECT 80.520 154.030 83.300 160.910 ;
        RECT 104.380 159.030 109.660 169.950 ;
        RECT 111.920 169.390 112.280 172.990 ;
        RECT 113.000 172.990 114.440 174.190 ;
        RECT 113.000 169.390 113.360 172.990 ;
        RECT 114.080 169.390 114.440 172.990 ;
        RECT 115.160 172.990 116.600 174.190 ;
        RECT 115.160 169.390 115.520 172.990 ;
        RECT 111.920 159.790 113.360 162.190 ;
        RECT 114.080 159.790 115.520 162.190 ;
        RECT 117.780 159.030 119.020 174.950 ;
        RECT 85.560 154.790 87.000 157.190 ;
        RECT 87.720 154.790 89.160 157.190 ;
        RECT 89.880 154.790 91.320 157.190 ;
        RECT 92.040 154.790 93.480 157.190 ;
        RECT 94.200 154.790 95.640 157.190 ;
        RECT 96.360 154.790 97.800 157.190 ;
        RECT 98.520 154.790 99.960 157.190 ;
        RECT 100.680 154.790 102.120 157.190 ;
        RECT 104.380 156.950 119.020 159.030 ;
        RECT 104.380 156.190 109.660 156.950 ;
        RECT 104.380 154.990 112.280 156.190 ;
        RECT 104.380 154.030 109.660 154.990 ;
        RECT 68.620 153.440 69.460 153.460 ;
        RECT 65.920 153.140 69.520 153.440 ;
        RECT 64.120 152.740 65.620 153.040 ;
        RECT 70.420 152.740 71.320 153.040 ;
        RECT 13.020 151.890 63.220 152.695 ;
        RECT 13.020 136.030 13.660 151.890 ;
        RECT 14.840 149.990 16.280 151.190 ;
        RECT 15.920 146.390 16.280 149.990 ;
        RECT 17.000 149.990 18.440 151.190 ;
        RECT 17.000 146.390 17.360 149.990 ;
        RECT 18.080 146.390 18.440 149.990 ;
        RECT 19.160 149.990 20.600 151.190 ;
        RECT 19.160 146.390 19.520 149.990 ;
        RECT 20.240 146.390 20.600 149.990 ;
        RECT 21.320 149.990 22.760 151.190 ;
        RECT 21.320 146.390 21.680 149.990 ;
        RECT 22.400 146.390 22.760 149.990 ;
        RECT 23.480 149.990 24.920 151.190 ;
        RECT 23.480 146.390 23.840 149.990 ;
        RECT 24.560 146.390 24.920 149.990 ;
        RECT 25.640 149.990 27.080 151.190 ;
        RECT 25.640 146.390 26.000 149.990 ;
        RECT 26.720 146.390 27.080 149.990 ;
        RECT 27.800 149.990 29.240 151.190 ;
        RECT 27.800 146.390 28.160 149.990 ;
        RECT 28.880 146.390 29.240 149.990 ;
        RECT 29.960 149.990 31.400 151.190 ;
        RECT 29.960 146.390 30.320 149.990 ;
        RECT 31.040 146.390 31.400 149.990 ;
        RECT 32.120 149.990 33.560 151.190 ;
        RECT 32.120 146.390 32.480 149.990 ;
        RECT 34.740 148.785 63.220 151.890 ;
        RECT 65.320 151.840 65.620 152.740 ;
        RECT 65.920 152.640 66.760 152.660 ;
        RECT 68.620 152.640 69.460 152.660 ;
        RECT 65.920 152.340 66.820 152.640 ;
        RECT 68.620 152.340 69.520 152.640 ;
        RECT 65.920 151.840 66.760 151.860 ;
        RECT 65.320 151.540 69.520 151.840 ;
        RECT 64.120 151.440 64.960 151.460 ;
        RECT 64.120 151.140 65.020 151.440 ;
        RECT 69.820 151.140 71.320 151.440 ;
        RECT 65.920 150.740 69.520 151.040 ;
        RECT 64.120 150.340 65.020 150.640 ;
        RECT 65.920 149.940 66.820 150.240 ;
        RECT 64.120 149.840 64.960 149.860 ;
        RECT 64.120 149.540 65.020 149.840 ;
        RECT 65.920 149.440 66.760 149.460 ;
        RECT 68.020 149.440 68.320 150.740 ;
        RECT 68.620 150.240 69.460 150.260 ;
        RECT 68.620 149.940 69.520 150.240 ;
        RECT 65.920 149.140 66.820 149.440 ;
        RECT 68.020 149.140 69.520 149.440 ;
        RECT 34.740 144.695 39.325 148.785 ;
        RECT 39.635 145.005 43.105 148.475 ;
        RECT 43.415 144.695 47.325 148.785 ;
        RECT 47.635 145.005 51.105 148.475 ;
        RECT 51.415 144.695 55.325 148.785 ;
        RECT 55.635 145.005 59.105 148.475 ;
        RECT 59.415 144.695 63.220 148.785 ;
        RECT 65.920 148.640 66.760 148.660 ;
        RECT 65.920 148.340 69.520 148.640 ;
        RECT 64.120 147.940 65.020 148.240 ;
        RECT 64.720 147.640 65.620 147.940 ;
        RECT 64.120 147.140 65.020 147.440 ;
        RECT 64.120 145.840 64.960 145.860 ;
        RECT 64.120 145.540 65.020 145.840 ;
        RECT 34.740 140.785 63.220 144.695 ;
        RECT 65.320 144.240 65.620 147.640 ;
        RECT 65.920 147.540 66.820 147.840 ;
        RECT 68.620 147.540 69.520 147.840 ;
        RECT 65.920 147.040 66.760 147.060 ;
        RECT 68.620 147.040 69.460 147.060 ;
        RECT 65.920 146.740 66.820 147.040 ;
        RECT 68.620 146.740 69.520 147.040 ;
        RECT 68.620 146.240 69.460 146.260 ;
        RECT 65.920 145.940 69.520 146.240 ;
        RECT 65.920 145.440 66.760 145.460 ;
        RECT 68.620 145.440 69.460 145.460 ;
        RECT 65.920 145.140 66.820 145.440 ;
        RECT 68.620 145.140 69.520 145.440 ;
        RECT 65.920 144.640 66.760 144.660 ;
        RECT 65.920 144.340 69.520 144.640 ;
        RECT 64.120 143.940 65.620 144.240 ;
        RECT 64.120 143.140 65.020 143.440 ;
        RECT 64.120 141.840 64.960 141.860 ;
        RECT 64.120 141.540 65.020 141.840 ;
        RECT 15.920 136.790 17.360 139.190 ;
        RECT 18.080 136.790 19.520 139.190 ;
        RECT 20.240 136.790 21.680 139.190 ;
        RECT 22.400 136.790 23.840 139.190 ;
        RECT 24.560 136.790 26.000 139.190 ;
        RECT 26.720 136.790 28.160 139.190 ;
        RECT 28.880 136.790 30.320 139.190 ;
        RECT 31.040 136.790 32.480 139.190 ;
        RECT 34.740 136.695 39.325 140.785 ;
        RECT 39.635 137.005 43.105 140.475 ;
        RECT 43.415 136.695 47.325 140.785 ;
        RECT 47.635 137.005 51.105 140.475 ;
        RECT 51.415 136.695 55.325 140.785 ;
        RECT 55.635 137.005 59.105 140.475 ;
        RECT 59.415 136.695 63.220 140.785 ;
        RECT 64.120 140.740 65.020 141.040 ;
        RECT 65.320 139.840 65.620 143.940 ;
        RECT 65.920 143.540 66.820 143.840 ;
        RECT 65.920 143.040 66.760 143.060 ;
        RECT 65.920 142.740 66.820 143.040 ;
        RECT 67.120 142.240 67.420 144.340 ;
        RECT 68.620 143.540 69.520 143.840 ;
        RECT 68.620 143.040 69.460 143.060 ;
        RECT 68.620 142.740 69.520 143.040 ;
        RECT 65.920 141.940 69.520 142.240 ;
        RECT 69.820 141.840 70.120 151.140 ;
        RECT 70.420 150.640 71.260 150.660 ;
        RECT 70.420 150.340 71.320 150.640 ;
        RECT 70.420 149.540 71.320 149.840 ;
        RECT 70.420 148.240 71.260 148.260 ;
        RECT 70.420 147.940 71.320 148.240 ;
        RECT 70.420 147.440 71.260 147.460 ;
        RECT 70.420 147.140 71.320 147.440 ;
        RECT 70.420 145.540 71.320 145.840 ;
        RECT 70.420 144.240 71.260 144.260 ;
        RECT 70.420 143.940 71.320 144.240 ;
        RECT 70.420 143.440 71.260 143.460 ;
        RECT 70.420 143.140 71.320 143.440 ;
        RECT 69.820 141.540 71.320 141.840 ;
        RECT 65.920 141.140 66.820 141.440 ;
        RECT 68.620 141.140 69.520 141.440 ;
        RECT 65.920 140.640 66.760 140.660 ;
        RECT 68.620 140.640 69.460 140.660 ;
        RECT 65.920 140.340 66.820 140.640 ;
        RECT 68.620 140.340 69.520 140.640 ;
        RECT 69.820 139.840 70.120 141.540 ;
        RECT 70.420 140.740 71.320 141.040 ;
        RECT 70.870 140.240 71.170 140.740 ;
        RECT 65.320 139.540 70.120 139.840 ;
        RECT 64.120 139.140 65.020 139.440 ;
        RECT 70.420 139.140 71.320 139.440 ;
        RECT 65.920 139.040 66.760 139.060 ;
        RECT 68.620 139.040 69.460 139.060 ;
        RECT 65.920 138.740 66.820 139.040 ;
        RECT 68.620 138.740 69.520 139.040 ;
        RECT 69.820 138.840 70.720 139.140 ;
        RECT 65.920 138.240 66.760 138.260 ;
        RECT 68.620 138.240 69.460 138.260 ;
        RECT 65.920 137.940 67.420 138.240 ;
        RECT 68.620 137.940 69.520 138.240 ;
        RECT 64.120 137.840 64.960 137.860 ;
        RECT 64.120 137.540 65.020 137.840 ;
        RECT 67.120 137.440 67.420 137.940 ;
        RECT 68.620 137.440 69.460 137.460 ;
        RECT 69.820 137.440 70.120 138.840 ;
        RECT 70.420 137.540 71.320 137.840 ;
        RECT 65.920 137.140 66.820 137.440 ;
        RECT 67.120 137.140 70.120 137.440 ;
        RECT 63.870 136.740 65.020 137.040 ;
        RECT 70.420 136.740 71.320 137.040 ;
        RECT 34.740 136.030 63.220 136.695 ;
        RECT 65.920 136.640 66.760 136.660 ;
        RECT 68.620 136.640 69.460 136.660 ;
        RECT 65.920 136.340 66.820 136.640 ;
        RECT 68.620 136.340 69.520 136.640 ;
        RECT 13.020 135.440 63.220 136.030 ;
        RECT 65.920 135.840 66.760 135.860 ;
        RECT 68.620 135.840 69.460 135.860 ;
        RECT 65.320 135.540 66.820 135.840 ;
        RECT 68.620 135.540 70.120 135.840 ;
        RECT 65.320 135.440 65.620 135.540 ;
        RECT 13.020 135.140 65.620 135.440 ;
        RECT 13.020 134.290 63.220 135.140 ;
        RECT 65.320 135.040 65.620 135.140 ;
        RECT 69.820 135.440 70.120 135.540 ;
        RECT 72.220 135.440 73.120 153.890 ;
        RECT 80.520 153.390 109.660 154.030 ;
        RECT 69.820 135.140 73.120 135.440 ;
        RECT 65.920 135.040 66.760 135.060 ;
        RECT 68.620 135.040 69.460 135.060 ;
        RECT 69.820 135.040 70.120 135.140 ;
        RECT 65.320 134.740 66.820 135.040 ;
        RECT 68.620 134.740 70.120 135.040 ;
        RECT 13.020 133.890 63.020 134.290 ;
        RECT 13.020 118.030 13.660 133.890 ;
        RECT 14.840 131.990 16.280 133.190 ;
        RECT 15.920 128.390 16.280 131.990 ;
        RECT 17.000 131.990 18.440 133.190 ;
        RECT 17.000 128.390 17.360 131.990 ;
        RECT 18.080 128.390 18.440 131.990 ;
        RECT 19.160 131.990 20.600 133.190 ;
        RECT 19.160 128.390 19.520 131.990 ;
        RECT 20.240 128.390 20.600 131.990 ;
        RECT 21.320 131.990 22.760 133.190 ;
        RECT 21.320 128.390 21.680 131.990 ;
        RECT 22.400 128.390 22.760 131.990 ;
        RECT 23.480 131.990 24.920 133.190 ;
        RECT 23.480 128.390 23.840 131.990 ;
        RECT 24.560 128.390 24.920 131.990 ;
        RECT 25.640 131.990 27.080 133.190 ;
        RECT 25.640 128.390 26.000 131.990 ;
        RECT 26.720 128.390 27.080 131.990 ;
        RECT 27.800 131.990 29.240 133.190 ;
        RECT 27.800 128.390 28.160 131.990 ;
        RECT 28.880 128.390 29.240 131.990 ;
        RECT 29.960 131.990 31.400 133.190 ;
        RECT 29.960 128.390 30.320 131.990 ;
        RECT 31.040 128.390 31.400 131.990 ;
        RECT 32.120 131.990 33.560 133.190 ;
        RECT 32.120 128.390 32.480 131.990 ;
        RECT 15.920 118.790 17.360 121.190 ;
        RECT 18.080 118.790 19.520 121.190 ;
        RECT 20.240 118.790 21.680 121.190 ;
        RECT 22.400 118.790 23.840 121.190 ;
        RECT 24.560 118.790 26.000 121.190 ;
        RECT 26.720 118.790 28.160 121.190 ;
        RECT 28.880 118.790 30.320 121.190 ;
        RECT 31.040 118.790 32.480 121.190 ;
        RECT 34.740 118.030 37.660 133.890 ;
        RECT 38.840 131.990 40.280 133.190 ;
        RECT 39.920 128.390 40.280 131.990 ;
        RECT 41.000 131.990 42.440 133.190 ;
        RECT 41.000 128.390 41.360 131.990 ;
        RECT 42.080 128.390 42.440 131.990 ;
        RECT 43.160 131.990 44.600 133.190 ;
        RECT 43.160 128.390 43.520 131.990 ;
        RECT 44.240 128.390 44.600 131.990 ;
        RECT 45.320 131.990 46.760 133.190 ;
        RECT 45.320 128.390 45.680 131.990 ;
        RECT 46.400 128.390 46.760 131.990 ;
        RECT 47.480 131.990 48.920 133.190 ;
        RECT 47.480 128.390 47.840 131.990 ;
        RECT 48.560 128.390 48.920 131.990 ;
        RECT 49.640 131.990 51.080 133.190 ;
        RECT 49.640 128.390 50.000 131.990 ;
        RECT 50.720 128.390 51.080 131.990 ;
        RECT 51.800 131.990 53.240 133.190 ;
        RECT 51.800 128.390 52.160 131.990 ;
        RECT 52.880 128.390 53.240 131.990 ;
        RECT 53.960 131.990 55.400 133.190 ;
        RECT 53.960 128.390 54.320 131.990 ;
        RECT 55.040 128.390 55.400 131.990 ;
        RECT 56.120 131.990 57.560 133.190 ;
        RECT 56.120 128.390 56.480 131.990 ;
        RECT 58.740 124.370 60.920 133.890 ;
        RECT 69.670 133.840 69.970 134.740 ;
        RECT 72.220 134.290 73.120 135.140 ;
        RECT 77.020 141.030 109.660 153.390 ;
        RECT 111.920 151.390 112.280 154.990 ;
        RECT 113.000 154.990 114.440 156.190 ;
        RECT 113.000 151.390 113.360 154.990 ;
        RECT 114.080 151.390 114.440 154.990 ;
        RECT 115.160 154.990 116.600 156.190 ;
        RECT 115.160 151.390 115.520 154.990 ;
        RECT 111.920 141.790 113.360 144.190 ;
        RECT 114.080 141.790 115.520 144.190 ;
        RECT 117.780 141.030 119.020 156.950 ;
        RECT 77.020 139.890 119.020 141.030 ;
        RECT 77.020 136.390 105.020 139.890 ;
        RECT 65.080 132.890 66.040 133.530 ;
        RECT 77.020 132.890 85.520 136.390 ;
        RECT 61.880 131.930 63.480 132.330 ;
        RECT 61.240 130.730 61.560 131.930 ;
        RECT 62.520 131.130 64.120 131.530 ;
        RECT 64.440 130.730 64.760 131.930 ;
        RECT 61.880 130.330 63.480 130.730 ;
        RECT 61.880 127.130 63.480 127.530 ;
        RECT 61.240 125.930 61.560 127.130 ;
        RECT 62.520 126.330 64.120 126.730 ;
        RECT 64.440 125.930 64.760 127.130 ;
        RECT 61.880 125.530 63.480 125.930 ;
        RECT 65.080 124.370 85.520 132.890 ;
        RECT 58.740 121.890 85.520 124.370 ;
        RECT 39.920 118.790 41.360 121.190 ;
        RECT 42.080 118.790 43.520 121.190 ;
        RECT 44.240 118.790 45.680 121.190 ;
        RECT 46.400 118.790 47.840 121.190 ;
        RECT 48.560 118.790 50.000 121.190 ;
        RECT 50.720 118.790 52.160 121.190 ;
        RECT 52.880 118.790 54.320 121.190 ;
        RECT 55.040 118.790 56.480 121.190 ;
        RECT 58.740 118.030 59.520 121.890 ;
        RECT 13.020 117.390 59.520 118.030 ;
      LAYER met1 ;
        RECT 12.520 211.990 108.520 212.390 ;
        RECT 12.520 211.870 108.620 211.990 ;
        RECT 12.380 210.390 108.620 211.870 ;
        RECT 11.740 189.870 12.060 209.330 ;
        RECT 12.380 191.230 13.340 210.390 ;
        RECT 14.300 189.870 15.260 209.330 ;
        RECT 20.740 189.870 21.060 208.830 ;
        RECT 21.380 191.230 22.340 210.390 ;
        RECT 23.300 205.880 24.260 208.830 ;
        RECT 23.290 193.860 24.270 205.880 ;
        RECT 23.300 189.870 24.260 193.860 ;
        RECT 29.740 189.870 30.060 208.830 ;
        RECT 30.380 191.230 31.340 210.390 ;
        RECT 32.300 189.870 33.260 208.830 ;
        RECT 38.740 189.870 39.060 208.830 ;
        RECT 39.380 191.230 40.340 210.390 ;
        RECT 41.300 189.870 42.260 208.830 ;
        RECT 47.740 201.710 48.060 201.830 ;
        RECT 47.420 189.870 48.060 201.710 ;
        RECT 48.380 198.230 49.340 210.390 ;
        RECT 11.540 189.230 48.060 189.870 ;
        RECT 11.540 188.910 48.000 189.230 ;
        RECT 32.360 187.290 33.560 188.910 ;
        RECT 50.300 187.930 51.260 201.830 ;
        RECT 56.740 189.050 57.060 208.830 ;
        RECT 57.380 191.230 58.340 210.390 ;
        RECT 59.300 204.370 60.260 208.830 ;
        RECT 59.270 203.410 60.290 204.370 ;
        RECT 59.300 195.880 60.260 201.830 ;
        RECT 49.570 187.870 51.260 187.930 ;
        RECT 53.860 188.730 57.060 189.050 ;
        RECT 59.300 188.880 60.260 194.830 ;
        RECT 13.420 185.890 16.120 187.290 ;
        RECT 32.220 185.890 33.720 187.290 ;
        RECT 39.380 186.910 51.300 187.870 ;
        RECT 13.420 169.290 14.620 185.890 ;
        RECT 38.740 175.230 39.060 186.580 ;
        RECT 39.380 175.230 40.340 186.910 ;
        RECT 41.300 173.870 42.260 186.330 ;
        RECT 47.740 175.230 48.060 186.580 ;
        RECT 48.380 175.230 49.340 186.910 ;
        RECT 49.570 186.850 50.530 186.910 ;
        RECT 38.540 172.910 48.500 173.870 ;
        RECT 50.300 173.550 51.260 185.830 ;
        RECT 53.860 173.550 54.180 188.730 ;
        RECT 50.300 173.030 54.180 173.550 ;
        RECT 13.420 167.890 16.120 169.290 ;
        RECT 38.740 162.230 39.060 172.910 ;
        RECT 39.380 161.860 40.340 170.830 ;
        RECT 41.300 162.230 42.260 172.910 ;
        RECT 47.740 162.230 48.060 172.910 ;
        RECT 44.510 161.870 45.470 161.930 ;
        RECT 48.380 161.870 49.340 170.830 ;
        RECT 50.300 162.230 51.260 173.030 ;
        RECT 53.860 166.550 54.180 173.030 ;
        RECT 53.860 166.230 56.210 166.550 ;
        RECT 43.600 161.860 49.340 161.870 ;
        RECT 39.380 160.920 49.340 161.860 ;
        RECT 39.380 160.910 40.340 160.920 ;
        RECT 43.600 160.910 49.340 160.920 ;
        RECT 44.510 160.850 45.470 160.910 ;
        RECT 35.890 159.050 37.150 160.250 ;
        RECT 61.520 159.670 63.520 210.390 ;
        RECT 66.780 187.930 67.740 201.830 ;
        RECT 68.700 198.230 69.660 210.390 ;
        RECT 69.980 201.710 70.300 201.830 ;
        RECT 69.980 189.870 70.620 201.710 ;
        RECT 75.780 189.870 76.740 208.830 ;
        RECT 77.700 191.230 78.660 210.390 ;
        RECT 78.980 189.870 79.300 208.830 ;
        RECT 84.780 189.870 85.740 208.830 ;
        RECT 86.700 191.230 87.660 210.390 ;
        RECT 87.980 189.870 88.300 208.830 ;
        RECT 93.780 205.880 94.740 208.830 ;
        RECT 93.770 193.860 94.750 205.880 ;
        RECT 93.780 189.870 94.740 193.860 ;
        RECT 95.700 191.230 96.660 210.390 ;
        RECT 96.980 189.870 97.300 208.830 ;
        RECT 102.780 189.870 103.740 209.330 ;
        RECT 104.700 191.230 105.660 210.390 ;
        RECT 107.420 210.190 108.620 210.390 ;
        RECT 110.720 210.190 112.120 210.290 ;
        RECT 105.980 189.870 106.300 209.330 ;
        RECT 107.420 208.990 112.120 210.190 ;
        RECT 110.720 208.890 112.120 208.990 ;
        RECT 115.320 208.890 117.620 210.290 ;
        RECT 116.420 192.290 117.620 208.890 ;
        RECT 109.920 190.890 112.120 192.290 ;
        RECT 115.320 190.890 117.620 192.290 ;
        RECT 69.980 189.230 106.500 189.870 ;
        RECT 70.040 188.910 106.500 189.230 ;
        RECT 66.780 187.870 68.470 187.930 ;
        RECT 66.740 186.910 78.660 187.870 ;
        RECT 84.480 187.290 85.680 188.910 ;
        RECT 67.510 186.850 68.470 186.910 ;
        RECT 66.780 173.440 67.740 185.830 ;
        RECT 68.700 175.230 69.660 186.910 ;
        RECT 69.980 175.230 70.300 186.580 ;
        RECT 75.780 173.870 76.740 186.330 ;
        RECT 77.700 175.230 78.660 186.910 ;
        RECT 78.980 175.230 79.300 186.580 ;
        RECT 84.320 185.890 85.820 187.290 ;
        RECT 101.920 185.890 104.620 187.290 ;
        RECT 64.270 173.140 67.740 173.440 ;
        RECT 64.270 160.340 64.570 173.140 ;
        RECT 66.780 162.230 67.740 173.140 ;
        RECT 69.540 172.910 79.500 173.870 ;
        RECT 68.700 161.870 69.660 170.830 ;
        RECT 69.980 162.230 70.300 172.910 ;
        RECT 75.780 162.230 76.740 172.910 ;
        RECT 72.570 161.870 73.530 161.930 ;
        RECT 68.700 161.860 74.440 161.870 ;
        RECT 77.700 161.860 78.660 170.830 ;
        RECT 78.980 162.230 79.300 172.910 ;
        RECT 103.420 169.290 104.620 185.890 ;
        RECT 109.920 174.250 111.120 190.890 ;
        RECT 116.600 174.250 117.620 176.230 ;
        RECT 109.920 172.990 112.010 174.250 ;
        RECT 110.810 172.930 112.010 172.990 ;
        RECT 115.430 172.930 117.620 174.250 ;
        RECT 101.920 167.890 104.620 169.290 ;
        RECT 68.700 160.920 78.660 161.860 ;
        RECT 68.700 160.910 74.440 160.920 ;
        RECT 77.700 160.910 78.660 160.920 ;
        RECT 72.570 160.850 73.530 160.910 ;
        RECT 64.270 160.040 72.600 160.340 ;
        RECT 13.920 149.890 16.120 151.290 ;
        RECT 32.390 151.190 33.590 151.250 ;
        RECT 35.920 151.190 37.120 159.050 ;
        RECT 61.520 158.710 65.830 159.670 ;
        RECT 51.170 158.440 51.470 158.470 ;
        RECT 49.940 158.140 51.470 158.440 ;
        RECT 51.170 158.110 51.470 158.140 ;
        RECT 32.390 149.990 37.120 151.190 ;
        RECT 39.620 153.090 59.120 156.490 ;
        RECT 61.520 156.390 63.520 158.710 ;
        RECT 65.940 156.010 66.240 158.600 ;
        RECT 66.740 157.440 67.620 157.780 ;
        RECT 69.440 157.440 70.320 157.780 ;
        RECT 72.300 156.980 72.600 160.040 ;
        RECT 71.080 156.330 71.960 156.360 ;
        RECT 71.080 155.450 75.190 156.330 ;
        RECT 116.420 156.250 117.620 172.930 ;
        RECT 71.080 155.420 71.960 155.450 ;
        RECT 115.430 154.990 117.620 156.250 ;
        RECT 115.430 154.930 116.630 154.990 ;
        RECT 67.840 154.040 68.140 154.100 ;
        RECT 65.340 153.740 68.140 154.040 ;
        RECT 67.840 153.680 68.140 153.740 ;
        RECT 68.620 153.440 69.500 153.480 ;
        RECT 68.620 153.140 70.120 153.440 ;
        RECT 32.390 149.930 33.590 149.990 ;
        RECT 13.920 133.290 15.120 149.890 ;
        RECT 39.620 140.390 43.020 153.090 ;
        RECT 48.920 148.265 50.120 151.020 ;
        RECT 47.845 145.215 50.895 148.265 ;
        RECT 55.820 140.390 59.120 153.090 ;
        RECT 65.920 152.340 66.800 152.680 ;
        RECT 68.620 152.340 69.500 152.680 ;
        RECT 65.920 151.840 66.800 151.880 ;
        RECT 65.920 151.540 67.420 151.840 ;
        RECT 64.120 151.140 65.000 151.480 ;
        RECT 64.120 149.840 65.000 149.880 ;
        RECT 39.620 137.090 59.120 140.390 ;
        RECT 63.520 149.540 65.000 149.840 ;
        RECT 63.520 137.840 63.820 149.540 ;
        RECT 65.920 149.140 66.800 149.480 ;
        RECT 65.920 148.640 66.800 148.680 ;
        RECT 67.120 148.640 67.420 151.540 ;
        RECT 69.820 150.640 70.120 153.140 ;
        RECT 102.890 152.490 104.090 152.550 ;
        RECT 100.890 151.290 104.090 152.490 ;
        RECT 102.890 151.230 104.090 151.290 ;
        RECT 70.420 150.640 71.300 150.680 ;
        RECT 69.820 150.340 71.300 150.640 ;
        RECT 68.620 149.940 69.500 150.280 ;
        RECT 65.920 148.340 67.420 148.640 ;
        RECT 70.420 148.240 71.300 148.280 ;
        RECT 70.420 147.940 71.920 148.240 ;
        RECT 70.420 147.440 71.300 147.480 ;
        RECT 69.820 147.140 71.300 147.440 ;
        RECT 65.920 146.740 66.800 147.080 ;
        RECT 68.620 146.740 69.500 147.080 ;
        RECT 68.620 146.240 69.500 146.280 ;
        RECT 69.820 146.240 70.120 147.140 ;
        RECT 68.620 145.940 70.120 146.240 ;
        RECT 64.120 145.840 65.000 145.880 ;
        RECT 64.120 145.540 65.620 145.840 ;
        RECT 65.320 144.640 65.620 145.540 ;
        RECT 65.920 145.140 66.800 145.480 ;
        RECT 68.620 145.140 69.500 145.480 ;
        RECT 65.920 144.640 66.800 144.680 ;
        RECT 65.320 144.340 66.800 144.640 ;
        RECT 69.820 143.440 70.120 145.940 ;
        RECT 70.420 144.240 71.300 144.280 ;
        RECT 71.620 144.240 71.920 147.940 ;
        RECT 70.420 143.940 71.920 144.240 ;
        RECT 70.420 143.440 71.300 143.480 ;
        RECT 69.820 143.140 71.300 143.440 ;
        RECT 65.920 142.740 66.800 143.080 ;
        RECT 68.620 142.740 69.500 143.080 ;
        RECT 64.120 141.840 65.000 141.880 ;
        RECT 64.120 141.540 65.020 141.840 ;
        RECT 64.720 141.240 65.620 141.540 ;
        RECT 65.320 138.240 65.620 141.240 ;
        RECT 65.920 140.340 66.800 140.680 ;
        RECT 68.620 140.340 69.500 140.680 ;
        RECT 70.810 140.210 71.230 140.510 ;
        RECT 70.870 139.710 71.170 140.210 ;
        RECT 65.920 138.740 66.800 139.080 ;
        RECT 68.620 138.740 69.500 139.080 ;
        RECT 65.920 138.240 66.800 138.280 ;
        RECT 65.320 137.940 66.800 138.240 ;
        RECT 68.620 137.940 69.500 138.280 ;
        RECT 64.120 137.840 65.000 137.880 ;
        RECT 63.520 137.540 65.000 137.840 ;
        RECT 56.360 133.290 57.560 137.090 ;
        RECT 63.520 134.140 63.820 137.540 ;
        RECT 68.620 137.440 69.500 137.480 ;
        RECT 71.620 137.440 71.920 143.940 ;
        RECT 68.620 137.140 71.920 137.440 ;
        RECT 65.920 136.340 66.800 136.680 ;
        RECT 68.620 136.340 69.500 136.680 ;
        RECT 65.920 135.540 66.800 135.880 ;
        RECT 68.620 135.540 69.500 135.880 ;
        RECT 65.920 134.740 66.800 135.080 ;
        RECT 68.620 134.740 69.500 135.080 ;
        RECT 63.520 133.840 70.000 134.140 ;
        RECT 13.920 131.890 16.220 133.290 ;
        RECT 32.320 133.190 33.620 133.290 ;
        RECT 38.720 133.190 40.120 133.290 ;
        RECT 32.320 131.990 40.120 133.190 ;
        RECT 32.320 131.890 33.620 131.990 ;
        RECT 38.720 131.890 40.120 131.990 ;
        RECT 56.320 131.890 57.620 133.290 ;
        RECT 61.170 132.740 61.620 133.190 ;
        RECT 61.240 124.730 61.560 132.740 ;
        RECT 61.880 123.380 62.840 133.130 ;
        RECT 63.160 132.170 67.430 133.130 ;
        RECT 63.160 124.730 64.120 132.170 ;
        RECT 66.700 129.140 67.640 130.020 ;
        RECT 66.730 127.610 67.610 129.140 ;
      LAYER met2 ;
        RECT 59.300 204.370 60.260 204.400 ;
        RECT 59.300 203.410 64.145 204.370 ;
        RECT 59.300 203.380 60.260 203.410 ;
        RECT 53.495 195.910 60.290 196.870 ;
        RECT 53.420 188.790 60.620 189.990 ;
        RECT 63.620 189.600 108.120 190.290 ;
        RECT 63.620 189.090 108.130 189.600 ;
        RECT 38.740 186.550 39.060 188.595 ;
        RECT 53.420 186.550 54.620 188.790 ;
        RECT 38.710 186.230 39.090 186.550 ;
        RECT 47.710 186.230 54.620 186.550 ;
        RECT 53.420 164.790 54.620 186.230 ;
        RECT 63.620 186.550 64.820 189.090 ;
        RECT 78.980 186.550 79.300 188.595 ;
        RECT 63.620 186.230 70.330 186.550 ;
        RECT 78.950 186.230 79.330 186.550 ;
        RECT 63.620 185.890 64.820 186.230 ;
        RECT 106.920 176.200 108.130 189.090 ;
        RECT 106.920 175.190 117.650 176.200 ;
        RECT 107.110 175.180 117.650 175.190 ;
        RECT 55.860 166.550 56.180 166.580 ;
        RECT 55.860 166.230 57.225 166.550 ;
        RECT 55.860 166.200 56.180 166.230 ;
        RECT 36.170 164.490 63.170 164.790 ;
        RECT 35.920 160.250 37.120 160.280 ;
        RECT 35.920 159.050 43.965 160.250 ;
        RECT 35.920 159.020 37.120 159.050 ;
        RECT 52.680 158.440 52.960 158.475 ;
        RECT 51.140 158.140 52.970 158.440 ;
        RECT 52.680 158.105 52.960 158.140 ;
        RECT 53.420 150.990 54.620 164.490 ;
        RECT 64.840 159.670 65.800 159.700 ;
        RECT 64.840 158.710 67.645 159.670 ;
        RECT 64.840 158.680 65.800 158.710 ;
        RECT 66.740 157.440 67.620 157.780 ;
        RECT 69.440 157.440 70.320 157.780 ;
        RECT 65.910 156.040 66.270 156.340 ;
        RECT 69.440 156.305 71.990 156.330 ;
        RECT 65.940 154.540 66.240 156.040 ;
        RECT 69.420 155.475 71.990 156.305 ;
        RECT 69.440 155.450 71.990 155.475 ;
        RECT 65.940 154.240 72.170 154.540 ;
        RECT 65.370 154.040 65.670 154.070 ;
        RECT 61.370 153.930 65.670 154.040 ;
        RECT 48.890 149.790 54.620 150.990 ;
        RECT 61.240 153.740 65.670 153.930 ;
        RECT 61.240 133.190 61.560 153.740 ;
        RECT 65.370 153.710 65.670 153.740 ;
        RECT 65.920 152.340 66.800 152.680 ;
        RECT 68.620 152.340 69.500 152.680 ;
        RECT 64.120 151.440 65.000 151.480 ;
        RECT 64.120 151.140 65.620 151.440 ;
        RECT 65.320 148.240 65.620 151.140 ;
        RECT 68.620 149.940 69.500 150.280 ;
        RECT 65.920 149.140 66.800 149.480 ;
        RECT 70.420 148.240 71.300 148.280 ;
        RECT 65.320 147.940 71.300 148.240 ;
        RECT 65.920 146.740 66.800 147.080 ;
        RECT 68.620 146.740 69.500 147.080 ;
        RECT 65.920 145.140 66.800 145.480 ;
        RECT 68.620 145.140 69.500 145.480 ;
        RECT 65.920 142.740 66.800 143.080 ;
        RECT 68.620 142.740 69.500 143.080 ;
        RECT 65.920 140.340 66.800 140.680 ;
        RECT 68.620 140.340 69.500 140.680 ;
        RECT 71.870 140.040 72.170 154.240 ;
        RECT 100.920 152.490 102.120 152.520 ;
        RECT 98.875 151.290 102.120 152.490 ;
        RECT 100.920 151.260 102.120 151.290 ;
        RECT 70.840 139.740 72.170 140.040 ;
        RECT 65.920 138.740 66.800 139.080 ;
        RECT 68.620 138.740 69.500 139.080 ;
        RECT 68.620 137.940 69.500 138.280 ;
        RECT 65.920 136.340 66.800 136.680 ;
        RECT 68.620 136.340 69.500 136.680 ;
        RECT 65.920 135.540 66.800 135.880 ;
        RECT 68.620 135.540 69.500 135.880 ;
        RECT 65.920 134.740 66.800 135.080 ;
        RECT 68.620 134.740 69.500 135.080 ;
        RECT 61.170 132.740 61.620 133.190 ;
        RECT 66.440 133.130 67.400 133.160 ;
        RECT 66.440 132.170 70.345 133.130 ;
        RECT 66.440 132.140 67.400 132.170 ;
        RECT 66.730 131.815 67.610 131.840 ;
        RECT 66.710 130.985 67.630 131.815 ;
        RECT 66.730 129.110 67.610 130.985 ;
      LAYER met3 ;
        RECT 38.715 188.570 39.085 188.575 ;
        RECT 53.420 188.570 54.620 196.990 ;
        RECT 38.715 188.250 54.620 188.570 ;
        RECT 38.715 188.245 39.085 188.250 ;
        RECT 42.745 160.250 43.945 160.275 ;
        RECT 53.420 160.250 54.620 188.250 ;
        RECT 63.165 188.970 64.125 204.395 ;
        RECT 63.165 188.010 82.700 188.970 ;
        RECT 56.875 166.550 57.205 166.575 ;
        RECT 56.860 166.230 59.680 166.550 ;
        RECT 56.875 166.205 57.205 166.230 ;
        RECT 59.360 164.790 59.680 166.230 ;
        RECT 42.745 159.050 54.620 160.250 ;
        RECT 56.120 159.390 61.520 164.790 ;
        RECT 42.745 159.025 43.945 159.050 ;
        RECT 52.655 158.440 52.985 158.455 ;
        RECT 54.960 158.440 55.280 158.480 ;
        RECT 52.655 158.140 55.280 158.440 ;
        RECT 52.655 158.125 52.985 158.140 ;
        RECT 54.960 158.100 55.280 158.140 ;
        RECT 66.665 155.270 67.625 159.695 ;
        RECT 69.440 155.450 70.320 158.790 ;
        RECT 66.665 154.830 69.200 155.270 ;
        RECT 66.665 154.310 69.500 154.830 ;
        RECT 65.920 131.840 66.800 153.690 ;
        RECT 68.620 134.490 69.500 154.310 ;
        RECT 81.740 151.590 82.700 188.010 ;
        RECT 98.895 152.490 100.095 152.515 ;
        RECT 79.020 146.190 84.420 151.590 ;
        RECT 86.820 146.190 92.220 151.590 ;
        RECT 96.890 151.290 100.095 152.490 ;
        RECT 98.895 151.265 100.095 151.290 ;
        RECT 81.520 143.790 81.920 146.190 ;
        RECT 89.320 143.790 89.720 146.190 ;
        RECT 79.020 140.370 84.420 143.790 ;
        RECT 74.540 139.410 84.420 140.370 ;
        RECT 69.365 133.130 70.325 133.155 ;
        RECT 74.540 133.130 75.500 139.410 ;
        RECT 79.020 138.890 84.420 139.410 ;
        RECT 86.820 138.890 92.220 143.790 ;
        RECT 79.020 138.390 92.220 138.890 ;
        RECT 69.365 132.170 75.500 133.130 ;
        RECT 69.365 132.145 70.325 132.170 ;
        RECT 65.920 130.960 67.610 131.840 ;
      LAYER met4 ;
        RECT 56.120 159.390 61.520 164.790 ;
        RECT 54.955 158.440 55.285 158.455 ;
        RECT 57.570 158.440 57.870 159.390 ;
        RECT 54.955 158.140 57.870 158.440 ;
        RECT 54.955 158.125 55.285 158.140 ;
        RECT 79.020 146.190 84.420 151.590 ;
        RECT 86.820 150.490 92.220 151.590 ;
        RECT 96.915 150.490 98.115 152.495 ;
        RECT 86.820 149.290 98.115 150.490 ;
        RECT 86.820 146.190 92.220 149.290 ;
        RECT 81.520 143.790 81.920 146.190 ;
        RECT 89.320 143.790 89.720 146.190 ;
        RECT 79.020 138.890 84.420 143.790 ;
        RECT 86.820 138.890 92.220 143.790 ;
        RECT 79.020 138.390 92.220 138.890 ;
  END
END tt_um_jnw_wulffern
END LIBRARY

