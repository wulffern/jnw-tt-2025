** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TT_SKY130A/tt_um_jnw_wulffern.sch
.subckt tt_um_jnw_wulffern VDPWR VGND ui_in<7> ui_in<6> ui_in<5> ui_in<4> ui_in<3> ui_in<2> ui_in<1> ui_in<0>
+ uo_out<7> uo_out<6> uo_out<5> uo_out<4> uo_out<3> uo_out<2> uo_out<1> uo_out<0> uio_in<7> uio_in<6> uio_in<5> uio_in<4> uio_in<3> uio_in<2> uio_in<1> uio_in<0>
+ uio_out<7> uio_out<6> uio_out<5> uio_out<4> uio_out<3> uio_out<2> uio_out<1> uio_out<0> ena clk rst_n uio_oe<7> uio_oe<6> uio_oe<5> uio_oe<4> uio_oe<3> uio_oe<2> uio_oe<1> uio_oe<0>
*.ipin VDPWR
*.ipin VGND
*.ipin ui_in<7> ui_in<6> ui_in<5> ui_in<4> ui_in<3> ui_in<2> ui_in<1> ui_in<0>
*.opin uo_out<7> uo_out<6> uo_out<5> uo_out<4> uo_out<3> uo_out<2> uo_out<1> uo_out<0>
*.ipin uio_in<7> uio_in<6> uio_in<5> uio_in<4> uio_in<3> uio_in<2> uio_in<1> uio_in<0>
*.opin uio_out<7> uio_out<6> uio_out<5> uio_out<4> uio_out<3> uio_out<2> uio_out<1> uio_out<0>
*.ipin ena
*.ipin clk
*.ipin rst_n
*.opin uio_oe<7> uio_oe<6> uio_oe<5> uio_oe<4> uio_oe<3> uio_oe<2> uio_oe<1> uio_oe<0>
x1 VDPWR OUT06 RST VGND JNW_GR06
x2 VDPWR VGND net1 CLK_B JNW_GR07
x3 ui_in<0> RST VDPWR VGND JNWTR_BFX1_CV
x4 OUT06 uo_out<1> VDPWR VGND JNWTR_BFX1_CV
x5 net1 uo_out<0> VDPWR VGND JNWTR_BFX1_CV
x6 RST net2 VDPWR VGND JNWTR_IVX1_CV
x7 RST OUT06 uo_out<2> VDPWR VGND JNWTR_NRX1_CV
x8 VDPWR VGND JNWTR_TAPCELLB_CV
x9 TIE_L VDPWR VGND JNWTR_TIEL_CV
R1<7> TIE_L uio_oe<7> sky130_fd_pr__res_generic_m4 W=0.3 L=0.3 m=1
R1<6> TIE_L uio_oe<6> sky130_fd_pr__res_generic_m4 W=0.3 L=0.3 m=1
R1<5> TIE_L uio_oe<5> sky130_fd_pr__res_generic_m4 W=0.3 L=0.3 m=1
R1<4> TIE_L uio_oe<4> sky130_fd_pr__res_generic_m4 W=0.3 L=0.3 m=1
R1<3> TIE_L uio_oe<3> sky130_fd_pr__res_generic_m4 W=0.3 L=0.3 m=1
R1<2> TIE_L uio_oe<2> sky130_fd_pr__res_generic_m4 W=0.3 L=0.3 m=1
R1<1> TIE_L uio_oe<1> sky130_fd_pr__res_generic_m4 W=0.3 L=0.3 m=1
R1<0> TIE_L uio_oe<0> sky130_fd_pr__res_generic_m4 W=0.3 L=0.3 m=1
x10 clk CLK_B VDPWR VGND JNWTR_BFX1_CV
.ends

* expanding   symbol:  JNW_GR06_SKY130A/JNW_GR06.sym # of pins=4
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_GR06_SKY130A/JNW_GR06.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_GR06_SKY130A/JNW_GR06.sch
.subckt JNW_GR06 VDD OUT reset VSS
*.ipin VDD
*.ipin VSS
*.opin OUT
*.ipin reset
x1 VDD CAP VSS temp_affected_current
x5 net2 net1 VSS JNWTR_RPPO4
x6 net1 VSS VSS JNWTR_RPPO4
x7 VDD net2 VSS JNWTR_RPPO4
x3 VDD CAP net1 OUT VSS OTA
x2 CAP VSS JNWTR_CAPX1
x4 CAP reset VSS VSS JNWATR_NCH_2C1F2
.ends


* expanding   symbol:  JNW_GR07_SKY130A/JNW_GR07.sym # of pins=4
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_GR07_SKY130A/JNW_GR07.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_GR07_SKY130A/JNW_GR07.sch
.subckt JNW_GR07 VDD VSS PWM CLK
*.ipin VDD
*.opin PWM
*.ipin VSS
*.ipin CLK
x3 V_OUT_OPAMP Buffer VDD VSS JNWTR_BFX1_CV
x5 Buffer CLK VDD PWM net3 VDD VSS JNWTR_DFRNQNX1_CV
x2<1> V_C PWM VSS VSS JNWATR_NCH_2C1F2
x2<0> V_C PWM VSS VSS JNWATR_NCH_2C1F2
x8 VSS V_REF VSS JNWTR_RPPO4
x9 V_REF net2 VSS JNWTR_RPPO4
x10 net2 net1 VSS JNWTR_RPPO4
x6 net1 VDD VSS JNWTR_RPPO4
x7 V_C VSS JNWTR_CAPX4
x4 VDD V_C V_REF V_OUT_OPAMP VSS amplifier_rev2
x11 VDD V_C VSS temp_to_current_rev2
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_BFX1_CV.sym # of pins=4
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_BFX1_CV.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_BFX1_CV.sch
.subckt JNWTR_BFX1_CV A Y AVDD AVSS
*.ipin A
*.opin Y
*.ipin AVDD
*.ipin AVSS
XMN0 AVSS A B AVSS JNWTR_NCHDL
XMN1 Y B AVSS AVSS JNWTR_NCHDL
XMP0 AVDD A B AVDD JNWTR_PCHDL
XMP1 Y B AVDD AVDD JNWTR_PCHDL
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_IVX1_CV.sym # of pins=4
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_IVX1_CV.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_IVX1_CV.sch
.subckt JNWTR_IVX1_CV A Y AVDD AVSS
*.ipin A
*.opin Y
*.ipin AVDD
*.ipin AVSS
XMN0 Y A AVSS AVSS JNWTR_NCHDL
XMP0 Y A AVDD AVDD JNWTR_PCHDL
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_NRX1_CV.sym # of pins=5
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_NRX1_CV.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_NRX1_CV.sch
.subckt JNWTR_NRX1_CV A B Y AVDD AVSS
*.iopin A
*.iopin B
*.iopin Y
*.iopin AVDD
*.iopin AVSS
XMN0 Y A AVSS AVSS JNWTR_NCHDL
XMN1 AVSS B Y AVSS JNWTR_NCHDL
XMP0 N1 A AVDD AVDD JNWTR_PCHDL
XMP1 Y B N1 AVDD JNWTR_PCHDL
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_TAPCELLB_CV.sym # of pins=2
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_TAPCELLB_CV.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_TAPCELLB_CV.sch
.subckt JNWTR_TAPCELLB_CV AVDD AVSS
*.iopin AVDD
*.iopin AVSS
XMN1 AVSS AVSS AVSS AVSS JNWTR_NCHDL
XMP1 AVDD AVDD AVDD AVDD JNWTR_PCHDL
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_TIEL_CV.sym # of pins=3
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_TIEL_CV.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_TIEL_CV.sch
.subckt JNWTR_TIEL_CV Y AVDD AVSS
*.iopin Y
*.iopin AVDD
*.iopin AVSS
XMN0 Y A AVSS AVSS JNWTR_NCHDL
XMP0 A A AVDD AVDD JNWTR_PCHDL
.ends


* expanding   symbol:  JNW_GR06_SKY130A/temp_affected_current.sym # of pins=3
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_GR06_SKY130A/temp_affected_current.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_GR06_SKY130A/temp_affected_current.sch
.subckt temp_affected_current VDD OUT VSS
*.ipin VDD
*.ipin VSS
*.opin OUT
x1 RIGHT_SIDE GATE VDD VDD JNWATR_PCH_4C5F0
x2 LEFT_SIDE GATE VDD VDD JNWATR_PCH_4C5F0
x3 VDD RIGHT_SIDE LEFT_SIDE GATE VSS OTA
XxQ1 VSS VSS LEFT_SIDE sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1 mult=1
XxQ2 VSS VSS VR sky130_fd_pr__pnp_05v5_W3p40L3p40 m=8 mult=8
x8 VDD GATE JNWTR_CAPX1
x4 net1 GATE VDD VDD JNWATR_PCH_4C5F0
x10<9> net2 net2 VDD VDD JNWATR_PCH_4C5F0
x10<8> net2 net2 VDD VDD JNWATR_PCH_4C5F0
x10<7> net2 net2 VDD VDD JNWATR_PCH_4C5F0
x10<6> net2 net2 VDD VDD JNWATR_PCH_4C5F0
x10<5> net2 net2 VDD VDD JNWATR_PCH_4C5F0
x10<4> net2 net2 VDD VDD JNWATR_PCH_4C5F0
x10<3> net2 net2 VDD VDD JNWATR_PCH_4C5F0
x10<2> net2 net2 VDD VDD JNWATR_PCH_4C5F0
x10<1> net2 net2 VDD VDD JNWATR_PCH_4C5F0
x10<0> net2 net2 VDD VDD JNWATR_PCH_4C5F0
x9 OUT net2 VDD VDD JNWATR_PCH_4C5F0
x5<9> net1 net1 VSS VSS JNWATR_NCH_4C5F0
x5<8> net1 net1 VSS VSS JNWATR_NCH_4C5F0
x5<7> net1 net1 VSS VSS JNWATR_NCH_4C5F0
x5<6> net1 net1 VSS VSS JNWATR_NCH_4C5F0
x5<5> net1 net1 VSS VSS JNWATR_NCH_4C5F0
x5<4> net1 net1 VSS VSS JNWATR_NCH_4C5F0
x5<3> net1 net1 VSS VSS JNWATR_NCH_4C5F0
x5<2> net1 net1 VSS VSS JNWATR_NCH_4C5F0
x5<1> net1 net1 VSS VSS JNWATR_NCH_4C5F0
x5<0> net1 net1 VSS VSS JNWATR_NCH_4C5F0
x6 net2 net1 VSS VSS JNWATR_NCH_4C5F0
x7 net3 VR VSS JNWTR_RPPO8
x10 RIGHT_SIDE net3 VSS JNWTR_RPPO4
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO4.sym # of pins=3
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO4.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO4.sch
.subckt JNWTR_RPPO4 N P B
*.iopin P
*.iopin N
*.iopin B
XXA1 N P B JNWTR_RES4
.ends


* expanding   symbol:  JNW_GR06_SKY130A/OTA.sym # of pins=5
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_GR06_SKY130A/OTA.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_GR06_SKY130A/OTA.sch
.subckt OTA VDD IN+ IN- OUT VSS
*.ipin IN+
*.ipin IN-
*.ipin VDD
*.ipin VSS
*.opin OUT
xd3<3> GATE IN+ OTA_SPLIT OTA_SPLIT JNWATR_PCH_4C5F0
xd3<2> GATE IN+ OTA_SPLIT OTA_SPLIT JNWATR_PCH_4C5F0
xd3<1> GATE IN+ OTA_SPLIT OTA_SPLIT JNWATR_PCH_4C5F0
xd3<0> GATE IN+ OTA_SPLIT OTA_SPLIT JNWATR_PCH_4C5F0
xe3<3> OUT IN- OTA_SPLIT OTA_SPLIT JNWATR_PCH_4C5F0
xe3<2> OUT IN- OTA_SPLIT OTA_SPLIT JNWATR_PCH_4C5F0
xe3<1> OUT IN- OTA_SPLIT OTA_SPLIT JNWATR_PCH_4C5F0
xe3<0> OUT IN- OTA_SPLIT OTA_SPLIT JNWATR_PCH_4C5F0
xa4b OTA_SPLIT IB_GATE VDD VDD JNWATR_PCH_4C5F0
xa4a IB_GATE IB_GATE VDD VDD JNWATR_PCH_4C5F0
xa1 VSS AFTER_RESISTOR2 VSS JNWTR_RPPO16
xa2 AFTER_RESISTOR2 AFTER_RESISTOR1 VSS JNWTR_RPPO16
xa3 AFTER_RESISTOR1 IB_GATE VSS JNWTR_RPPO16
xd2 GATE GATE VSS VSS JNWATR_NCH_4C5F0
xe2 OUT GATE VSS VSS JNWATR_NCH_4C5F0
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_CAPX1.sym # of pins=2
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sch
.subckt JNWTR_CAPX1 A B
*.iopin A
*.iopin B
XC1 B A sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_2C1F2.sym # of pins=4
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_2C1F2.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_2C1F2.sch
.subckt JNWATR_NCH_2C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.22 W=1.92 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_DFRNQNX1_CV.sym # of pins=7
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_DFRNQNX1_CV.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_DFRNQNX1_CV.sch
.subckt JNWTR_DFRNQNX1_CV D CK RN Q QN AVDD AVSS
*.iopin D
*.iopin CK
*.iopin RN
*.iopin Q
*.iopin QN
*.iopin AVDD
*.iopin AVSS
XXA0 AVDD AVSS JNWTR_TAPCELLB_CV
XXA1 CK RN CKN AVDD AVSS JNWTR_NDX1_CV
XXA2 CKN CKB AVDD AVSS JNWTR_IVX1_CV
XXA3 D CKN CKB A0 AVDD AVSS JNWTR_IVTRIX1_CV
XXA4 A1 CKB CKN A0 AVDD AVSS JNWTR_IVTRIX1_CV
XXA5 A0 A1 AVDD AVSS JNWTR_IVX1_CV
XXA6 A1 CKB CKN QN AVDD AVSS JNWTR_IVTRIX1_CV
XXA7 Q CKN CKB RN QN AVDD AVSS JNWTR_NDTRIX1_CV
XXA8 QN Q AVDD AVSS JNWTR_IVX1_CV
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_CAPX4.sym # of pins=2
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX4.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX4.sch
.subckt JNWTR_CAPX4 A B
*.iopin A
*.iopin B
XXA1 A B JNWTR_CAPX1
XXA2 A B JNWTR_CAPX1
XXB1 A B JNWTR_CAPX1
XXB2 A B JNWTR_CAPX1
.ends


* expanding   symbol:  JNW_GR07_SKY130A/amplifier_rev2.sym # of pins=5
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_GR07_SKY130A/amplifier_rev2.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_GR07_SKY130A/amplifier_rev2.sch
.subckt amplifier_rev2 VDD VINP VINN VOUT VSS
*.ipin VINP
*.ipin VINN
*.ipin VDD
*.ipin VSS
*.opin VOUT
x1<1> OTA_CM_gate OTA_CM_gate VSS VSS JNWATR_NCH_4C5F0
x1<0> OTA_CM_gate OTA_CM_gate VSS VSS JNWATR_NCH_4C5F0
x2<1> VOUT OTA_CM_gate VSS VSS JNWATR_NCH_4C5F0
x2<0> VOUT OTA_CM_gate VSS VSS JNWATR_NCH_4C5F0
x3<1> OTA_CM_gate VINP OTA_VDD OTA_VDD JNWATR_PCH_4C5F0
x3<0> OTA_CM_gate VINP OTA_VDD OTA_VDD JNWATR_PCH_4C5F0
x4<1> VOUT VINN OTA_VDD OTA_VDD JNWATR_PCH_4C5F0
x4<0> VOUT VINN OTA_VDD OTA_VDD JNWATR_PCH_4C5F0
x5 OTA_VDD IB_gate VDD VDD JNWATR_PCH_4C5F0
x6<11> IB_gate IB_gate VDD VDD JNWATR_PCH_4C5F0
x6<10> IB_gate IB_gate VDD VDD JNWATR_PCH_4C5F0
x6<9> IB_gate IB_gate VDD VDD JNWATR_PCH_4C5F0
x6<8> IB_gate IB_gate VDD VDD JNWATR_PCH_4C5F0
x6<7> IB_gate IB_gate VDD VDD JNWATR_PCH_4C5F0
x6<6> IB_gate IB_gate VDD VDD JNWATR_PCH_4C5F0
x6<5> IB_gate IB_gate VDD VDD JNWATR_PCH_4C5F0
x6<4> IB_gate IB_gate VDD VDD JNWATR_PCH_4C5F0
x6<3> IB_gate IB_gate VDD VDD JNWATR_PCH_4C5F0
x6<2> IB_gate IB_gate VDD VDD JNWATR_PCH_4C5F0
x6<1> IB_gate IB_gate VDD VDD JNWATR_PCH_4C5F0
x6<0> IB_gate IB_gate VDD VDD JNWATR_PCH_4C5F0
x4 VSS net1 VSS JNWTR_RPPO16
x1 net1 IB_gate VSS JNWTR_RPPO16
.ends


* expanding   symbol:  JNW_GR07_SKY130A/temp_to_current_rev2.sym # of pins=3
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_GR07_SKY130A/temp_to_current_rev2.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_GR07_SKY130A/temp_to_current_rev2.sch
.subckt temp_to_current_rev2 VDD I_OUT VSS
*.ipin VDD
*.opin I_OUT
*.ipin VSS
x VINP VOUT VDD VDD JNWATR_PCH_4C5F0
x3 VINN VOUT VDD VDD JNWATR_PCH_4C5F0
XQ1 VSS VSS VINN sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1 mult=1
XQ2 VSS VSS V_diode sky130_fd_pr__pnp_05v5_W3p40L3p40 m=8 mult=8
x5 I_OUT VOUT VDD VDD JNWATR_PCH_4C5F0
x2 VOUT VSS JNWTR_CAPX1
x4 net1 VINP VSS JNWTR_RPPO16
x6 net2 net1 VSS JNWTR_RPPO16
x7 V_diode net2 VSS JNWTR_RPPO16
x1 VDD VINP VINN VOUT VSS amplifier_rev2
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_NCHDL.sym # of pins=4
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_NCHDL.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_NCHDL.sch
.subckt JNWTR_NCHDL D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.16 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_PCHDL.sym # of pins=4
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_PCHDL.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_PCHDL.sch
.subckt JNWTR_PCHDL D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.16 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym # of pins=4
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sch
.subckt JNWATR_PCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym # of pins=4
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sch
.subckt JNWATR_NCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO8.sym # of pins=3
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO8.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO8.sch
.subckt JNWTR_RPPO8 N P B
*.iopin P
*.iopin N
*.iopin B
XXA1 N P B JNWTR_RES8
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES4.sym # of pins=3
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_RES4.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_RES4.sch
.subckt JNWTR_RES4 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 INT_1 INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_2 INT_2 INT_1 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_3 P INT_2 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO16.sym # of pins=3
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO16.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO16.sch
.subckt JNWTR_RPPO16 N P B
*.iopin P
*.iopin N
*.iopin B
XXA1 N P B JNWTR_RES16
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_NDX1_CV.sym # of pins=5
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_NDX1_CV.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_NDX1_CV.sch
.subckt JNWTR_NDX1_CV A B Y AVDD AVSS
*.iopin A
*.iopin B
*.iopin Y
*.iopin AVDD
*.iopin AVSS
XMN0 N1 A AVSS AVSS JNWTR_NCHDL
XMN1 Y B N1 AVSS JNWTR_NCHDL
XMP0 Y A AVDD AVDD JNWTR_PCHDL
XMP1 AVDD B Y AVDD JNWTR_PCHDL
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_IVTRIX1_CV.sym # of pins=6
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_IVTRIX1_CV.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_IVTRIX1_CV.sch
.subckt JNWTR_IVTRIX1_CV A C CN Y AVDD AVSS
*.iopin A
*.iopin C
*.iopin CN
*.iopin Y
*.iopin AVDD
*.iopin AVSS
XMN0 N1 A AVSS AVSS JNWTR_NCHDL
XMN1 Y C N1 AVSS JNWTR_NCHDL
XMP0 N2 A AVDD AVDD JNWTR_PCHDL
XMP1 Y CN N2 AVDD JNWTR_PCHDL
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_NDTRIX1_CV.sym # of pins=7
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_NDTRIX1_CV.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_NDTRIX1_CV.sch
.subckt JNWTR_NDTRIX1_CV A C CN RN Y AVDD AVSS
*.iopin A
*.iopin C
*.iopin CN
*.iopin RN
*.iopin Y
*.iopin AVDD
*.iopin AVSS
XMN2 N1 RN AVSS AVSS JNWTR_NCHDL
XMN0 N2 A N1 AVSS JNWTR_NCHDL
XMN1 Y C N2 AVSS JNWTR_NCHDL
XMP2 AVDD RN N2 AVDD JNWTR_PCHDL
XMP0 N2 A AVDD AVDD JNWTR_PCHDL
XMP1 Y CN N2 AVDD JNWTR_PCHDL
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES8.sym # of pins=3
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_RES8.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_RES8.sch
.subckt JNWTR_RES8 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 INT_1 INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_2 INT_2 INT_1 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_3 INT_3 INT_2 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_4 INT_4 INT_3 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_5 INT_5 INT_4 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_6 INT_6 INT_5 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_7 P INT_6 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES16.sym # of pins=3
** sym_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_RES16.sym
** sch_path: /Users/wulff/pro/jnw-tt-2025/ip/jnw_tt_sky130a/design/JNW_TR_SKY130A/JNWTR_RES16.sch
.subckt JNWTR_RES16 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 INT_1 INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_2 INT_2 INT_1 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_3 INT_3 INT_2 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_4 INT_4 INT_3 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_5 INT_5 INT_4 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_6 INT_6 INT_5 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_7 INT_7 INT_6 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_8 INT_8 INT_7 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_9 INT_9 INT_8 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_10 INT_10 INT_9 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_11 INT_11 INT_10 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_12 INT_12 INT_11 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_13 INT_13 INT_12 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_14 INT_14 INT_13 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_15 P INT_14 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends

.end
