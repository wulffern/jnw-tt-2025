magic
tech sky130A
magscale 1 2
timestamp 1755246527
<< locali >>
rect 4538 33530 4598 33536
rect 4538 33482 4544 33530
rect 4592 33482 4598 33530
rect 4538 33310 4598 33482
rect 3800 32996 3860 33096
rect 3800 32990 3974 32996
rect 3800 32942 3920 32990
rect 3968 32942 3974 32990
rect 3800 32936 3974 32942
rect 4364 32874 4486 32880
rect 4364 32826 4370 32874
rect 4418 32826 4486 32874
rect 4364 32820 4486 32826
rect 5110 32510 5174 32620
rect 5110 32458 5116 32510
rect 5168 32458 5174 32510
rect 5110 32452 5174 32458
rect 4072 32348 4178 32396
rect 4012 32336 4178 32348
rect 3812 32080 4048 32140
rect 3988 32076 4048 32080
rect 3988 32016 4584 32076
rect 3808 31472 3868 31836
rect 5065 31655 5132 31661
rect 5065 31600 5071 31655
rect 5126 31600 5132 31655
rect 5065 31467 5132 31600
rect 4042 31376 4392 31436
rect 3872 31306 3932 31360
rect 3830 31232 3932 31306
rect 3830 30900 3890 31232
rect 3830 30840 4062 30900
rect 4002 30796 4062 30840
rect 4880 30818 5126 30878
rect 4880 30796 4940 30818
rect 4002 30736 4396 30796
rect 4540 30736 4940 30796
rect 1944 27602 1966 27990
rect 2354 27988 2740 27990
rect 2354 27876 8833 27988
rect 2354 27712 4432 27876
rect 4596 27712 8833 27876
rect 2354 27602 8833 27712
rect 8447 27183 8833 27602
rect 21158 27236 21218 27388
rect 8447 26797 11035 27183
rect 4564 2686 5776 2692
rect 4564 2298 4570 2686
rect 4958 2298 5776 2686
rect 4564 2292 5776 2298
<< viali >>
rect 4544 33482 4592 33530
rect 3920 32942 3968 32990
rect 4370 32826 4418 32874
rect 5116 32458 5168 32510
rect 4012 32348 4072 32396
rect 3764 32080 3812 32140
rect 5071 31600 5126 31655
rect 3994 31376 4042 31436
rect 5126 30818 5174 30878
rect 3778 30496 3826 30556
rect 1966 27602 2354 27990
rect 4432 27712 4596 27876
rect 21158 27188 21218 27236
rect 4570 2298 4958 2686
<< metal1 >>
rect 4216 44704 4276 44710
rect 3914 44192 3974 44198
rect 2848 43876 2908 43882
rect 2578 43558 2638 43564
rect 2578 31442 2638 43498
rect 2848 32158 2908 43816
rect 3170 43692 3176 43752
rect 3236 43692 3242 43752
rect 2836 32140 2944 32158
rect 2836 32080 2850 32140
rect 2910 32080 2944 32140
rect 2836 32064 2944 32080
rect 2578 31436 2642 31442
rect 2578 31376 2582 31436
rect 2578 31370 2642 31376
rect 2578 31352 2638 31370
rect 3176 30556 3236 43692
rect 3914 32996 3974 44132
rect 4078 44020 4138 44026
rect 4078 33716 4138 43960
rect 4078 33650 4138 33656
rect 4216 33514 4276 44644
rect 11353 42620 11714 42626
rect 11714 42259 12176 42620
rect 11353 42253 11714 42259
rect 4538 34006 4598 34012
rect 4022 33454 4276 33514
rect 4364 33716 4424 33722
rect 3908 32990 3980 32996
rect 3908 32942 3920 32990
rect 3968 32942 3980 32990
rect 3908 32936 3980 32942
rect 4022 32824 4082 33454
rect 4012 32758 4082 32824
rect 4364 32874 4424 33656
rect 4538 33530 4598 33946
rect 4538 33482 4544 33530
rect 4592 33482 4598 33530
rect 4538 33470 4598 33482
rect 10052 34006 10112 34012
rect 4364 32826 4370 32874
rect 4418 32826 4424 32874
rect 4364 32814 4424 32826
rect 4012 32402 4072 32758
rect 5260 32600 5324 32606
rect 5260 32516 5324 32536
rect 5104 32510 5324 32516
rect 5104 32458 5116 32510
rect 5168 32458 5324 32510
rect 5104 32452 5324 32458
rect 9850 32600 9914 32606
rect 4000 32396 4084 32402
rect 4000 32348 4012 32396
rect 4072 32348 4084 32396
rect 4000 32342 4084 32348
rect 3758 32140 3818 32152
rect 3680 32080 3686 32140
rect 3746 32080 3764 32140
rect 3812 32080 3818 32140
rect 3758 32068 3818 32080
rect 5059 31655 5296 31661
rect 5059 31600 5071 31655
rect 5126 31600 5296 31655
rect 5059 31594 5296 31600
rect 5229 31506 5296 31594
rect 3988 31436 4048 31448
rect 5223 31439 5229 31506
rect 5296 31439 5302 31506
rect 3838 31376 3844 31436
rect 3904 31376 3994 31436
rect 4042 31376 4048 31436
rect 3988 31364 4048 31376
rect 5120 30878 5180 30890
rect 5756 30878 6000 32184
rect 6538 31568 6730 31770
rect 6532 31376 6538 31568
rect 6730 31376 6736 31568
rect 5120 30818 5126 30878
rect 5174 30818 5206 30878
rect 5266 30818 5272 30878
rect 5756 30818 5904 30878
rect 5964 30818 6000 30878
rect 5120 30806 5180 30818
rect 3772 30556 3832 30568
rect 3656 30496 3662 30556
rect 3722 30496 3778 30556
rect 3826 30496 3832 30556
rect 3176 30490 3236 30496
rect 3772 30484 3832 30496
rect 1232 27996 1632 28002
rect 1632 27990 2366 27996
rect 1632 27602 1966 27990
rect 2354 27602 2366 27990
rect 4112 27706 4118 27882
rect 4294 27876 4608 27882
rect 4294 27712 4432 27876
rect 4596 27712 4608 27876
rect 4294 27706 4608 27712
rect 1632 27596 2366 27602
rect 1232 27590 1632 27596
rect 5756 22194 6000 30818
rect 6538 22576 6730 31376
rect 9850 27260 9914 32536
rect 9850 27190 9914 27196
rect 10052 27112 10112 33946
rect 21146 27236 21230 27242
rect 21146 27188 21158 27236
rect 21218 27188 21230 27236
rect 21146 27182 21230 27188
rect 21158 27140 21218 27182
rect 10046 27052 10052 27112
rect 10112 27052 10118 27112
rect 21158 27074 21218 27080
rect 6538 22378 6730 22384
rect 31692 22576 31884 22582
rect 5756 21944 6000 21950
rect 6194 20760 6594 20766
rect 6594 20360 7574 20760
rect 6194 20354 6594 20360
rect 31692 19242 31884 22384
rect 30162 19050 31884 19242
rect 17618 10576 17624 10820
rect 17868 10576 18350 10820
rect 30162 7138 30354 19050
rect 29892 6946 30354 7138
rect 3584 2692 3984 2698
rect 3984 2686 4970 2692
rect 3984 2298 4570 2686
rect 4958 2298 4970 2686
rect 3984 2292 4970 2298
rect 3584 2286 3984 2292
<< via1 >>
rect 4216 44644 4276 44704
rect 3914 44132 3974 44192
rect 2848 43816 2908 43876
rect 2578 43498 2638 43558
rect 3176 43692 3236 43752
rect 2850 32080 2910 32140
rect 2582 31376 2642 31436
rect 4078 43960 4138 44020
rect 4078 33656 4138 33716
rect 11353 42259 11714 42620
rect 4538 33946 4598 34006
rect 4364 33656 4424 33716
rect 10052 33946 10112 34006
rect 5260 32536 5324 32600
rect 9850 32536 9914 32600
rect 3686 32080 3746 32140
rect 5229 31439 5296 31506
rect 3844 31376 3904 31436
rect 6538 31376 6730 31568
rect 5206 30818 5266 30878
rect 5904 30818 5964 30878
rect 3176 30496 3236 30556
rect 3662 30496 3722 30556
rect 1232 27596 1632 27996
rect 4118 27706 4294 27882
rect 9850 27196 9914 27260
rect 10052 27052 10112 27112
rect 21158 27080 21218 27140
rect 6538 22384 6730 22576
rect 31692 22384 31884 22576
rect 5756 21950 6000 22194
rect 6194 20360 6594 20760
rect 17624 10576 17868 10820
rect 3584 2292 3984 2692
<< metal2 >>
rect 4210 44644 4216 44704
rect 4276 44644 5510 44704
rect 5566 44644 5575 44704
rect 3908 44132 3914 44192
rect 3974 44190 28826 44192
rect 3974 44134 28768 44190
rect 28824 44134 28833 44190
rect 3974 44132 28826 44134
rect 18832 44020 18888 44027
rect 4072 43960 4078 44020
rect 4138 44018 18890 44020
rect 4138 43962 18832 44018
rect 18888 43962 18890 44018
rect 4138 43960 18890 43962
rect 18832 43953 18888 43960
rect 18280 43876 18336 43883
rect 2842 43816 2848 43876
rect 2908 43874 18338 43876
rect 2908 43818 18280 43874
rect 18336 43818 18338 43874
rect 2908 43816 18338 43818
rect 18280 43809 18336 43816
rect 3176 43752 3236 43758
rect 3236 43692 27654 43752
rect 27710 43692 27719 43752
rect 3176 43686 3236 43692
rect 2572 43498 2578 43558
rect 2638 43556 17786 43558
rect 2638 43500 17728 43556
rect 17784 43500 17793 43556
rect 2638 43498 17786 43500
rect 697 42616 11353 42620
rect 692 42615 11353 42616
rect 692 42611 4663 42615
rect 692 42221 697 42611
rect 1087 42449 4663 42611
rect 4829 42449 11353 42615
rect 1087 42259 11353 42449
rect 11714 42259 11720 42620
rect 1087 42221 1272 42259
rect 692 42216 1272 42221
rect 697 42212 1087 42216
rect 4532 33946 4538 34006
rect 4598 33946 10052 34006
rect 10112 33946 10118 34006
rect 4072 33656 4078 33716
rect 4138 33656 4364 33716
rect 4424 33656 4430 33716
rect 5254 32536 5260 32600
rect 5324 32536 9850 32600
rect 9914 32536 9920 32600
rect 3686 32140 3746 32146
rect 2844 32080 2850 32140
rect 2910 32080 3686 32140
rect 3686 32074 3746 32080
rect 6538 31568 6730 31574
rect 5229 31506 5296 31512
rect 3844 31436 3904 31442
rect 2576 31376 2582 31436
rect 2642 31376 3844 31436
rect 5296 31439 6538 31506
rect 5229 31433 5296 31439
rect 3844 31370 3904 31376
rect 6538 31370 6730 31376
rect 5206 30878 5266 30884
rect 5266 30818 5904 30878
rect 5964 30818 5970 30878
rect 5206 30812 5266 30818
rect 3662 30556 3722 30562
rect 3170 30496 3176 30556
rect 3236 30496 3662 30556
rect 3662 30490 3722 30496
rect 4118 28311 4294 28316
rect 4114 28145 4123 28311
rect 4289 28145 4298 28311
rect 805 27996 1195 28000
rect 800 27991 1232 27996
rect 800 27601 805 27991
rect 1195 27601 1232 27991
rect 800 27596 1232 27601
rect 1632 27596 1638 27996
rect 4118 27882 4294 28145
rect 4118 27700 4294 27706
rect 805 27592 1195 27596
rect 9844 27196 9850 27260
rect 9914 27196 20608 27260
rect 10052 27112 10112 27118
rect 10112 27052 20226 27112
rect 21152 27080 21158 27140
rect 21218 27080 21224 27140
rect 10052 27046 10112 27052
rect 20166 26408 20226 27052
rect 21158 26408 21218 27080
rect 20166 26348 21218 26408
rect 6532 22384 6538 22576
rect 6730 22384 31692 22576
rect 31884 22384 31890 22576
rect 5750 21950 5756 22194
rect 6000 22189 17249 22194
rect 6000 21955 17010 22189
rect 17244 21955 17253 22189
rect 6000 21950 17249 21955
rect 911 20760 1301 20764
rect 906 20755 6194 20760
rect 906 20365 911 20755
rect 1301 20365 6194 20755
rect 906 20360 6194 20365
rect 6594 20360 6600 20760
rect 911 20356 1301 20360
rect 17624 10820 17868 10826
rect 17001 10576 17010 10820
rect 17244 10576 17624 10820
rect 17624 10570 17868 10576
rect 2571 2692 2961 2696
rect 2566 2687 3584 2692
rect 2566 2297 2571 2687
rect 2961 2297 3584 2687
rect 2566 2292 3584 2297
rect 3984 2292 3990 2692
rect 2571 2288 2961 2292
<< via2 >>
rect 5510 44644 5566 44704
rect 28768 44134 28824 44190
rect 18832 43962 18888 44018
rect 18280 43818 18336 43874
rect 27654 43692 27710 43752
rect 17728 43500 17784 43556
rect 697 42221 1087 42611
rect 4663 42449 4829 42615
rect 4123 28145 4289 28311
rect 805 27601 1195 27991
rect 17010 21955 17244 22189
rect 911 20365 1301 20755
rect 17010 10576 17244 10820
rect 2571 2297 2961 2687
<< metal3 >>
rect 28758 44840 28764 44904
rect 28828 44840 28834 44904
rect 17718 44742 17724 44806
rect 17788 44742 17794 44806
rect 5505 44704 5571 44709
rect 6212 44704 6218 44706
rect 5505 44644 5510 44704
rect 5566 44644 6218 44704
rect 5505 44639 5571 44644
rect 6212 44642 6218 44644
rect 6282 44642 6288 44706
rect 17726 43561 17786 44742
rect 18270 44728 18276 44792
rect 18340 44728 18346 44792
rect 18822 44744 18828 44808
rect 18892 44744 18898 44808
rect 27650 44800 27714 44806
rect 18278 43879 18338 44728
rect 18830 44023 18890 44744
rect 27650 44730 27714 44736
rect 18827 44018 18893 44023
rect 18827 43962 18832 44018
rect 18888 43962 18893 44018
rect 18827 43957 18893 43962
rect 18275 43874 18341 43879
rect 18275 43818 18280 43874
rect 18336 43818 18341 43874
rect 18275 43813 18341 43818
rect 27652 43757 27712 44730
rect 28766 44195 28826 44840
rect 28763 44190 28829 44195
rect 28763 44134 28768 44190
rect 28824 44134 28829 44190
rect 28763 44129 28829 44134
rect 27649 43752 27715 43757
rect 27649 43692 27654 43752
rect 27710 43692 27715 43752
rect 27649 43687 27715 43692
rect 17723 43556 17789 43561
rect 17723 43500 17728 43556
rect 17784 43500 17789 43556
rect 17723 43495 17789 43500
rect 196 42616 608 42626
rect 196 42615 1092 42616
rect 196 42217 201 42615
rect 599 42611 1092 42615
rect 599 42221 697 42611
rect 1087 42221 1092 42611
rect 599 42217 1092 42221
rect 196 42216 1092 42217
rect 4658 42615 4834 42620
rect 4658 42449 4663 42615
rect 4829 42449 4834 42615
rect 196 42204 608 42216
rect 788 28683 1274 28742
rect 788 28285 801 28683
rect 1199 28285 1274 28683
rect 788 28276 1274 28285
rect 4118 28311 4294 32854
rect 4658 30396 4834 42449
rect 800 27991 1200 28276
rect 4118 28145 4123 28311
rect 4289 28145 4294 28311
rect 4118 28140 4294 28145
rect 800 27601 805 27991
rect 1195 27601 1200 27991
rect 800 27596 1200 27601
rect 17005 22189 17249 22194
rect 17005 21955 17010 22189
rect 17244 21955 17249 22189
rect 186 20760 672 20796
rect 186 20759 1306 20760
rect 186 20361 201 20759
rect 599 20755 1306 20759
rect 599 20365 911 20755
rect 1301 20365 1306 20755
rect 599 20361 1306 20365
rect 186 20360 1306 20361
rect 186 20330 672 20360
rect 17005 10820 17249 21955
rect 17005 10576 17010 10820
rect 17244 10576 17249 10820
rect 17005 10571 17249 10576
rect 748 2692 1234 2742
rect 748 2691 2966 2692
rect 748 2293 801 2691
rect 1199 2687 2966 2691
rect 1199 2297 2571 2687
rect 2961 2297 2966 2687
rect 1199 2293 2966 2297
rect 748 2292 2966 2293
rect 748 2276 1234 2292
<< via3 >>
rect 28764 44840 28828 44904
rect 17724 44742 17788 44806
rect 6218 44642 6282 44706
rect 18276 44728 18340 44792
rect 18828 44744 18892 44808
rect 27650 44736 27714 44800
rect 201 42217 599 42615
rect 801 28285 1199 28683
rect 201 20361 599 20759
rect 801 2293 1199 2691
<< metal4 >>
rect 6134 44868 6194 45152
rect 6134 44780 6194 44808
rect 6686 44874 6746 45152
rect 6686 44780 6746 44814
rect 7238 44876 7298 45152
rect 7238 44780 7298 44816
rect 7790 44878 7850 45152
rect 7790 44780 7850 44818
rect 8342 44876 8402 45152
rect 8342 44780 8402 44816
rect 8894 44870 8954 45152
rect 8894 44780 8954 44810
rect 9446 44884 9506 45152
rect 9446 44780 9506 44824
rect 9998 44914 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 9998 44871 10060 44914
rect 9998 44780 10060 44809
rect 17726 44807 17786 45152
rect 6134 44720 10060 44780
rect 17723 44806 17789 44807
rect 17723 44742 17724 44806
rect 17788 44742 17789 44806
rect 18278 44793 18338 45152
rect 18830 44809 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 45036 27722 45152
rect 27662 44970 27748 45036
rect 18827 44808 18893 44809
rect 17723 44741 17789 44742
rect 18275 44792 18341 44793
rect 18275 44728 18276 44792
rect 18340 44728 18341 44792
rect 18827 44744 18828 44808
rect 18892 44744 18893 44808
rect 18827 44743 18893 44744
rect 27622 44800 27770 44970
rect 28214 44952 28274 45152
rect 28766 44905 28826 45152
rect 29318 44952 29378 45152
rect 28763 44904 28829 44905
rect 28763 44840 28764 44904
rect 28828 44840 28829 44904
rect 28763 44839 28829 44840
rect 18275 44727 18341 44728
rect 27622 44736 27650 44800
rect 27714 44736 27770 44800
rect 27622 44726 27770 44736
rect 6142 44706 6384 44720
rect 6142 44642 6218 44706
rect 6282 44642 6384 44706
rect 6142 44618 6384 44642
rect 200 42615 600 44152
rect 200 42217 201 42615
rect 599 42217 600 42615
rect 200 20759 600 42217
rect 200 20361 201 20759
rect 599 20361 600 20759
rect 200 1000 600 20361
rect 800 28683 1200 44152
rect 800 28285 801 28683
rect 1199 28285 1200 28683
rect 800 2691 1200 28285
rect 800 2293 801 2691
rect 1199 2293 1200 2691
rect 800 1000 1200 2293
<< rmetal4 >>
rect 6134 44808 6194 44868
rect 6686 44814 6746 44874
rect 7238 44816 7298 44876
rect 7790 44818 7850 44878
rect 8342 44816 8402 44876
rect 8894 44810 8954 44870
rect 9446 44824 9506 44884
rect 9998 44809 10060 44871
use JNW_GR06  JNW_GR06_0 ../JNW_GR06_SKY130A
timestamp 1755246527
transform 1 0 904 0 1 3794
box -788 -2348 31548 17886
use JNW_GR07  JNW_GR07_0 ../JNW_GR07_SKY130A
timestamp 1755246527
transform 1 0 6300 0 1 31458
box 4000 -8000 25800 11000
use JNWTR_BFX1_CV  JNWTR_BFX1_CV_0 ../JNW_TR_SKY130A
timestamp 1755246527
transform 1 0 3488 0 1 30366
box -150 -120 2130 600
use JNWTR_BFX1_CV  JNWTR_BFX1_CV_1
timestamp 1755246527
transform 1 0 3488 0 1 32926
box -150 -120 2130 600
use JNWTR_BFX1_CV  JNWTR_BFX1_CV_2
timestamp 1755246527
transform 1 0 3488 0 1 31646
box -150 -120 2130 600
use JNWTR_BFX1_CV  JNWTR_BFX1_CV_3
timestamp 1755246527
transform 1 0 3488 0 1 32446
box -150 -120 2130 600
use JNWTR_IVX1_CV  JNWTR_IVX1_CV_0 ../JNW_TR_SKY130A
timestamp 1755246527
transform 1 0 3488 0 1 30846
box -150 -120 2130 440
use JNWTR_NRX1_CV  JNWTR_NRX1_CV_0 ../JNW_TR_SKY130A
timestamp 1755246527
transform 1 0 3488 0 1 31166
box -150 -120 2130 600
use JNWTR_TAPCELLB_CV  JNWTR_TAPCELLB_CV_0 ../JNW_TR_SKY130A
timestamp 1755246527
transform 1 0 3488 0 1 30046
box -150 -120 2130 440
use JNWTR_TIEL_CV  JNWTR_TIEL_CV_0 ../JNW_TR_SKY130A
timestamp 1755246527
transform 1 0 3488 0 1 32126
box -150 -120 2130 440
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal2 5148 44644 5208 44704 0 FreeSans 640 0 0 0 TIE_L
flabel metal2 6255 31439 6330 31506 0 FreeSans 640 0 0 0 OUT06
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
