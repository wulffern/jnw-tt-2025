MACRO tt_um_jnw_wulffern
  CLASS BLOCK ;
  FOREIGN tt_um_jnw_wulffern ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 10.020 204.890 17.620 210.170 ;
        RECT 19.020 204.390 26.620 209.670 ;
        RECT 28.020 204.390 35.620 209.670 ;
        RECT 37.020 204.390 44.620 209.670 ;
        RECT 55.020 204.390 62.620 209.670 ;
        RECT 73.420 204.390 81.020 209.670 ;
        RECT 82.420 204.390 90.020 209.670 ;
        RECT 91.420 204.390 99.020 209.670 ;
        RECT 100.420 204.890 108.020 210.170 ;
        RECT 10.020 197.390 17.620 202.670 ;
        RECT 19.020 197.390 26.620 202.670 ;
        RECT 28.020 197.390 35.620 202.670 ;
        RECT 37.020 197.390 44.620 202.670 ;
        RECT 46.020 197.390 53.620 202.670 ;
        RECT 55.020 197.390 62.620 202.670 ;
        RECT 64.420 197.390 72.020 202.670 ;
        RECT 73.420 197.390 81.020 202.670 ;
        RECT 82.420 197.390 90.020 202.670 ;
        RECT 91.420 197.390 99.020 202.670 ;
        RECT 100.420 197.390 108.020 202.670 ;
      LAYER pwell ;
        RECT 110.840 195.790 116.600 210.190 ;
      LAYER nwell ;
        RECT 10.020 190.390 17.620 195.670 ;
        RECT 19.020 190.390 26.620 195.670 ;
        RECT 28.020 190.390 35.620 195.670 ;
        RECT 37.020 190.390 44.620 195.670 ;
        RECT 55.020 190.390 62.620 195.670 ;
        RECT 73.420 190.390 81.020 195.670 ;
        RECT 82.420 190.390 90.020 195.670 ;
        RECT 91.420 190.390 99.020 195.670 ;
        RECT 100.420 190.390 108.020 195.670 ;
      LAYER pwell ;
        RECT 14.840 172.790 33.560 187.190 ;
      LAYER nwell ;
        RECT 37.020 181.890 44.620 187.170 ;
        RECT 46.020 181.390 53.620 186.670 ;
        RECT 64.420 181.390 72.020 186.670 ;
        RECT 73.420 181.890 81.020 187.170 ;
        RECT 37.020 174.390 44.620 179.670 ;
        RECT 46.020 174.390 53.620 179.670 ;
        RECT 64.420 174.390 72.020 179.670 ;
        RECT 73.420 174.390 81.020 179.670 ;
      LAYER pwell ;
        RECT 84.480 172.790 103.200 187.190 ;
        RECT 110.840 177.790 116.600 192.190 ;
        RECT 14.840 154.790 33.560 169.190 ;
        RECT 37.020 161.390 44.620 171.670 ;
        RECT 46.020 161.390 53.620 171.670 ;
        RECT 64.420 161.390 72.020 171.670 ;
        RECT 73.420 161.390 81.020 171.670 ;
        RECT 38.020 157.325 44.720 158.090 ;
        RECT 38.020 152.155 38.785 157.325 ;
        RECT 43.955 152.155 44.720 157.325 ;
        RECT 38.020 151.390 44.720 152.155 ;
        RECT 46.020 157.325 52.720 158.090 ;
        RECT 46.020 152.155 46.785 157.325 ;
        RECT 51.955 152.155 52.720 157.325 ;
        RECT 46.020 151.390 52.720 152.155 ;
        RECT 54.020 157.325 60.720 158.090 ;
        RECT 54.020 152.155 54.785 157.325 ;
        RECT 59.955 152.155 60.720 157.325 ;
      LAYER nwell ;
        RECT 62.820 155.790 68.520 159.390 ;
      LAYER pwell ;
        RECT 68.520 155.790 74.220 159.390 ;
        RECT 84.480 154.790 103.200 169.190 ;
        RECT 110.840 159.790 116.600 174.190 ;
        RECT 54.020 151.390 60.720 152.155 ;
        RECT 14.840 136.790 33.560 151.190 ;
        RECT 38.020 149.325 44.720 150.090 ;
        RECT 38.020 144.155 38.785 149.325 ;
        RECT 43.955 144.155 44.720 149.325 ;
        RECT 38.020 143.390 44.720 144.155 ;
        RECT 46.020 149.325 52.720 150.090 ;
        RECT 46.020 144.155 46.785 149.325 ;
        RECT 51.955 144.155 52.720 149.325 ;
        RECT 46.020 143.390 52.720 144.155 ;
        RECT 54.020 149.325 60.720 150.090 ;
        RECT 54.020 144.155 54.785 149.325 ;
        RECT 59.955 144.155 60.720 149.325 ;
        RECT 54.020 143.390 60.720 144.155 ;
        RECT 38.020 141.325 44.720 142.090 ;
        RECT 38.020 136.155 38.785 141.325 ;
        RECT 43.955 136.155 44.720 141.325 ;
        RECT 38.020 135.390 44.720 136.155 ;
        RECT 46.020 141.325 52.720 142.090 ;
        RECT 46.020 136.155 46.785 141.325 ;
        RECT 51.955 136.155 52.720 141.325 ;
        RECT 46.020 135.390 52.720 136.155 ;
        RECT 54.020 141.325 60.720 142.090 ;
        RECT 54.020 136.155 54.785 141.325 ;
        RECT 59.955 136.155 60.720 141.325 ;
        RECT 54.020 135.390 60.720 136.155 ;
        RECT 62.020 133.970 67.720 154.290 ;
        RECT 59.520 133.890 67.720 133.970 ;
      LAYER nwell ;
        RECT 67.720 133.890 73.420 154.290 ;
      LAYER pwell ;
        RECT 110.840 141.790 116.600 156.190 ;
        RECT 14.840 118.790 33.560 133.190 ;
        RECT 38.840 118.790 57.560 133.190 ;
        RECT 59.520 123.890 66.480 133.890 ;
      LAYER nwell ;
        RECT 73.740 96.610 81.340 100.770 ;
        RECT 73.720 95.490 81.340 96.610 ;
      LAYER pwell ;
        RECT 62.580 90.720 70.180 94.850 ;
      LAYER nwell ;
        RECT 73.720 92.620 81.320 95.490 ;
        RECT 73.720 91.330 81.360 92.620 ;
      LAYER pwell ;
        RECT 62.570 89.570 70.180 90.720 ;
        RECT 62.570 86.720 70.170 89.570 ;
      LAYER nwell ;
        RECT 73.760 88.460 81.360 91.330 ;
        RECT 73.720 87.340 81.360 88.460 ;
      LAYER pwell ;
        RECT 62.570 85.440 70.200 86.720 ;
        RECT 62.600 82.590 70.200 85.440 ;
      LAYER nwell ;
        RECT 73.720 84.460 81.320 87.340 ;
      LAYER pwell ;
        RECT 92.300 85.830 98.060 100.230 ;
        RECT 102.970 85.910 108.730 100.310 ;
        RECT 113.560 85.990 119.320 100.390 ;
      LAYER nwell ;
        RECT 73.720 83.180 81.340 84.460 ;
      LAYER pwell ;
        RECT 62.590 81.440 70.200 82.590 ;
        RECT 62.590 78.600 70.190 81.440 ;
      LAYER nwell ;
        RECT 73.740 80.300 81.340 83.180 ;
        RECT 73.720 79.180 81.340 80.300 ;
      LAYER pwell ;
        RECT 62.590 77.310 70.200 78.600 ;
        RECT 62.600 74.470 70.200 77.310 ;
      LAYER nwell ;
        RECT 73.720 76.170 81.320 79.180 ;
        RECT 73.720 75.020 81.340 76.170 ;
      LAYER pwell ;
        RECT 62.590 73.320 70.200 74.470 ;
        RECT 6.390 57.060 25.110 71.460 ;
        RECT 62.590 70.460 70.190 73.320 ;
      LAYER nwell ;
        RECT 73.740 72.010 81.340 75.020 ;
        RECT 73.740 70.890 81.350 72.010 ;
        RECT 33.330 64.190 40.930 69.210 ;
      LAYER pwell ;
        RECT 62.590 69.190 70.220 70.460 ;
        RECT 62.620 66.330 70.220 69.190 ;
      LAYER nwell ;
        RECT 73.750 67.880 81.350 70.890 ;
      LAYER pwell ;
        RECT 62.610 65.180 70.220 66.330 ;
      LAYER nwell ;
        RECT 73.730 66.730 81.350 67.880 ;
        RECT 33.330 63.930 40.950 64.190 ;
        RECT 33.350 58.910 40.950 63.930 ;
      LAYER pwell ;
        RECT 62.610 62.340 70.210 65.180 ;
      LAYER nwell ;
        RECT 73.730 63.720 81.330 66.730 ;
        RECT 73.730 62.600 81.350 63.720 ;
      LAYER pwell ;
        RECT 62.610 61.050 70.220 62.340 ;
        RECT 6.290 39.470 25.010 53.870 ;
      LAYER nwell ;
        RECT 28.580 48.840 36.180 57.140 ;
        RECT 38.490 48.880 46.090 57.180 ;
        RECT 54.110 53.620 61.710 58.900 ;
      LAYER pwell ;
        RECT 62.620 58.210 70.220 61.050 ;
      LAYER nwell ;
        RECT 73.750 58.440 81.350 62.600 ;
        RECT 83.100 58.440 90.700 63.720 ;
      LAYER pwell ;
        RECT 62.610 57.060 70.220 58.210 ;
        RECT 62.610 52.930 70.210 57.060 ;
        RECT 73.680 52.920 81.280 58.200 ;
        RECT 108.740 53.520 127.460 67.920 ;
      LAYER nwell ;
        RECT 135.680 60.650 143.280 65.670 ;
        RECT 135.680 60.390 143.300 60.650 ;
        RECT 135.700 55.370 143.300 60.390 ;
        RECT 28.570 47.750 36.180 48.840 ;
        RECT 38.480 47.790 46.090 48.880 ;
        RECT 28.570 39.450 36.170 47.750 ;
        RECT 38.480 39.490 46.080 47.790 ;
        RECT 59.760 39.170 67.360 43.290 ;
        RECT 59.760 38.010 67.370 39.170 ;
      LAYER pwell ;
        RECT 6.230 22.000 24.950 36.400 ;
        RECT 28.580 31.690 36.180 36.970 ;
        RECT 38.500 31.680 46.100 36.960 ;
      LAYER nwell ;
        RECT 59.770 33.890 67.370 38.010 ;
      LAYER pwell ;
        RECT 72.490 34.720 78.250 49.120 ;
        RECT 82.260 34.640 92.340 49.040 ;
        RECT 108.640 35.930 127.360 50.330 ;
      LAYER nwell ;
        RECT 130.930 45.300 138.530 53.600 ;
        RECT 140.840 45.340 148.440 53.640 ;
        RECT 130.920 44.210 138.530 45.300 ;
        RECT 140.830 44.250 148.440 45.340 ;
        RECT 130.920 35.910 138.520 44.210 ;
        RECT 140.830 35.950 148.430 44.250 ;
      LAYER pwell ;
        RECT 65.070 31.965 71.770 32.730 ;
        RECT 65.070 26.795 65.835 31.965 ;
        RECT 71.005 26.795 71.770 31.965 ;
        RECT 48.290 25.285 54.990 26.050 ;
        RECT 65.070 26.030 71.770 26.795 ;
        RECT 71.790 31.965 78.490 32.730 ;
        RECT 71.790 26.795 72.555 31.965 ;
        RECT 77.725 26.795 78.490 31.965 ;
        RECT 71.790 26.030 78.490 26.795 ;
        RECT 78.570 31.955 85.270 32.720 ;
        RECT 78.570 26.785 79.335 31.955 ;
        RECT 84.505 26.785 85.270 31.955 ;
        RECT 78.570 26.020 85.270 26.785 ;
        RECT 85.310 31.945 92.010 32.710 ;
        RECT 85.310 26.775 86.075 31.945 ;
        RECT 91.245 26.775 92.010 31.945 ;
        RECT 85.310 26.010 92.010 26.775 ;
        RECT 48.290 20.115 49.055 25.285 ;
        RECT 54.225 20.115 54.990 25.285 ;
        RECT 48.290 19.350 54.990 20.115 ;
        RECT 65.070 25.065 71.770 25.830 ;
        RECT 65.070 19.895 65.835 25.065 ;
        RECT 71.005 19.895 71.770 25.065 ;
        RECT 65.070 19.130 71.770 19.895 ;
        RECT 71.810 25.065 78.510 25.830 ;
        RECT 71.810 19.895 72.575 25.065 ;
        RECT 77.745 19.895 78.510 25.065 ;
        RECT 71.810 19.130 78.510 19.895 ;
        RECT 78.560 25.065 85.260 25.830 ;
        RECT 78.560 19.895 79.325 25.065 ;
        RECT 84.495 19.895 85.260 25.065 ;
        RECT 78.560 19.130 85.260 19.895 ;
        RECT 85.300 25.065 92.000 25.830 ;
        RECT 85.300 19.895 86.065 25.065 ;
        RECT 91.235 19.895 92.000 25.065 ;
        RECT 95.160 21.510 102.120 26.790 ;
        RECT 85.300 19.130 92.000 19.895 ;
        RECT 108.580 18.460 127.300 32.860 ;
        RECT 130.930 28.150 138.530 33.430 ;
        RECT 140.850 28.140 148.450 33.420 ;
      LAYER li1 ;
        RECT 10.520 210.870 107.520 211.890 ;
        RECT 109.020 210.950 119.020 211.890 ;
        RECT 10.460 209.910 107.580 210.870 ;
        RECT 10.460 190.870 11.420 209.910 ;
        RECT 12.380 208.930 14.620 209.330 ;
        RECT 11.740 206.930 12.060 208.130 ;
        RECT 13.020 207.330 15.260 207.730 ;
        RECT 15.580 206.930 15.900 208.130 ;
        RECT 12.380 205.730 14.620 206.130 ;
        RECT 12.380 201.430 14.620 201.830 ;
        RECT 11.740 199.430 12.060 200.630 ;
        RECT 13.020 199.830 15.260 200.230 ;
        RECT 15.580 199.430 15.900 200.630 ;
        RECT 12.380 198.230 14.620 198.630 ;
        RECT 12.380 194.430 14.620 194.830 ;
        RECT 11.740 192.430 12.060 193.630 ;
        RECT 13.020 192.830 15.260 193.230 ;
        RECT 15.580 192.430 15.900 193.630 ;
        RECT 12.380 191.230 14.620 191.630 ;
        RECT 16.220 190.870 20.420 209.910 ;
        RECT 21.380 208.430 23.620 208.830 ;
        RECT 20.740 206.430 21.060 207.630 ;
        RECT 22.020 206.830 24.260 207.230 ;
        RECT 24.580 206.430 24.900 207.630 ;
        RECT 21.380 205.230 23.620 205.630 ;
        RECT 21.380 201.430 23.620 201.830 ;
        RECT 20.740 199.430 21.060 200.630 ;
        RECT 22.020 199.830 24.260 200.230 ;
        RECT 24.580 199.430 24.900 200.630 ;
        RECT 21.380 198.230 23.620 198.630 ;
        RECT 21.380 194.430 23.620 194.830 ;
        RECT 20.740 192.430 21.060 193.630 ;
        RECT 22.020 192.830 24.260 193.230 ;
        RECT 24.580 192.430 24.900 193.630 ;
        RECT 21.380 191.230 23.620 191.630 ;
        RECT 25.220 190.870 29.420 209.910 ;
        RECT 30.380 208.430 32.620 208.830 ;
        RECT 29.740 206.430 30.060 207.630 ;
        RECT 31.020 206.830 33.260 207.230 ;
        RECT 33.580 206.430 33.900 207.630 ;
        RECT 30.380 205.230 32.620 205.630 ;
        RECT 30.380 201.430 32.620 201.830 ;
        RECT 29.740 199.430 30.060 200.630 ;
        RECT 31.020 199.830 33.260 200.230 ;
        RECT 33.580 199.430 33.900 200.630 ;
        RECT 30.380 198.230 32.620 198.630 ;
        RECT 30.380 194.430 32.620 194.830 ;
        RECT 29.740 192.430 30.060 193.630 ;
        RECT 31.020 192.830 33.260 193.230 ;
        RECT 33.580 192.430 33.900 193.630 ;
        RECT 30.380 191.230 32.620 191.630 ;
        RECT 34.220 190.870 38.420 209.910 ;
        RECT 39.380 208.430 41.620 208.830 ;
        RECT 38.740 206.430 39.060 207.630 ;
        RECT 40.020 206.830 42.260 207.230 ;
        RECT 42.580 206.430 42.900 207.630 ;
        RECT 39.380 205.230 41.620 205.630 ;
        RECT 43.220 202.410 56.420 209.910 ;
        RECT 57.380 208.430 59.620 208.830 ;
        RECT 56.740 206.430 57.060 207.630 ;
        RECT 58.020 206.830 60.260 207.230 ;
        RECT 60.580 206.430 60.900 207.630 ;
        RECT 57.380 205.230 59.620 205.630 ;
        RECT 39.380 201.430 41.620 201.830 ;
        RECT 38.740 199.430 39.060 200.630 ;
        RECT 40.020 199.830 42.260 200.230 ;
        RECT 42.580 199.430 42.900 200.630 ;
        RECT 39.380 198.230 41.620 198.630 ;
        RECT 43.220 197.870 47.420 202.410 ;
        RECT 48.380 201.430 50.620 201.830 ;
        RECT 47.740 199.430 48.060 200.630 ;
        RECT 49.020 199.830 51.260 200.230 ;
        RECT 51.580 199.430 51.900 200.630 ;
        RECT 48.380 198.230 50.620 198.630 ;
        RECT 52.220 197.870 56.420 202.410 ;
        RECT 61.220 202.410 74.820 209.910 ;
        RECT 76.420 208.430 78.660 208.830 ;
        RECT 75.140 206.430 75.460 207.630 ;
        RECT 75.780 206.830 78.020 207.230 ;
        RECT 78.980 206.430 79.300 207.630 ;
        RECT 76.420 205.230 78.660 205.630 ;
        RECT 57.380 201.430 59.620 201.830 ;
        RECT 56.740 199.430 57.060 200.630 ;
        RECT 58.020 199.830 60.260 200.230 ;
        RECT 60.580 199.430 60.900 200.630 ;
        RECT 57.380 198.230 59.620 198.630 ;
        RECT 39.380 194.430 41.620 194.830 ;
        RECT 38.740 192.430 39.060 193.630 ;
        RECT 40.020 192.830 42.260 193.230 ;
        RECT 42.580 192.430 42.900 193.630 ;
        RECT 39.380 191.230 41.620 191.630 ;
        RECT 43.220 190.870 56.420 197.870 ;
        RECT 61.220 197.870 65.820 202.410 ;
        RECT 67.420 201.430 69.660 201.830 ;
        RECT 66.140 199.430 66.460 200.630 ;
        RECT 66.780 199.830 69.020 200.230 ;
        RECT 69.980 199.430 70.300 200.630 ;
        RECT 67.420 198.230 69.660 198.630 ;
        RECT 70.620 197.870 74.820 202.410 ;
        RECT 76.420 201.430 78.660 201.830 ;
        RECT 75.140 199.430 75.460 200.630 ;
        RECT 75.780 199.830 78.020 200.230 ;
        RECT 78.980 199.430 79.300 200.630 ;
        RECT 76.420 198.230 78.660 198.630 ;
        RECT 57.380 194.430 59.620 194.830 ;
        RECT 56.740 192.430 57.060 193.630 ;
        RECT 58.020 192.830 60.260 193.230 ;
        RECT 60.580 192.430 60.900 193.630 ;
        RECT 57.380 191.230 59.620 191.630 ;
        RECT 61.220 190.870 74.820 197.870 ;
        RECT 76.420 194.430 78.660 194.830 ;
        RECT 75.140 192.430 75.460 193.630 ;
        RECT 75.780 192.830 78.020 193.230 ;
        RECT 78.980 192.430 79.300 193.630 ;
        RECT 76.420 191.230 78.660 191.630 ;
        RECT 79.620 190.870 83.820 209.910 ;
        RECT 85.420 208.430 87.660 208.830 ;
        RECT 84.140 206.430 84.460 207.630 ;
        RECT 84.780 206.830 87.020 207.230 ;
        RECT 87.980 206.430 88.300 207.630 ;
        RECT 85.420 205.230 87.660 205.630 ;
        RECT 85.420 201.430 87.660 201.830 ;
        RECT 84.140 199.430 84.460 200.630 ;
        RECT 84.780 199.830 87.020 200.230 ;
        RECT 87.980 199.430 88.300 200.630 ;
        RECT 85.420 198.230 87.660 198.630 ;
        RECT 85.420 194.430 87.660 194.830 ;
        RECT 84.140 192.430 84.460 193.630 ;
        RECT 84.780 192.830 87.020 193.230 ;
        RECT 87.980 192.430 88.300 193.630 ;
        RECT 85.420 191.230 87.660 191.630 ;
        RECT 88.620 190.870 92.820 209.910 ;
        RECT 94.420 208.430 96.660 208.830 ;
        RECT 93.140 206.430 93.460 207.630 ;
        RECT 93.780 206.830 96.020 207.230 ;
        RECT 96.980 206.430 97.300 207.630 ;
        RECT 94.420 205.230 96.660 205.630 ;
        RECT 94.420 201.430 96.660 201.830 ;
        RECT 93.140 199.430 93.460 200.630 ;
        RECT 93.780 199.830 96.020 200.230 ;
        RECT 96.980 199.430 97.300 200.630 ;
        RECT 94.420 198.230 96.660 198.630 ;
        RECT 94.420 194.430 96.660 194.830 ;
        RECT 93.140 192.430 93.460 193.630 ;
        RECT 93.780 192.830 96.020 193.230 ;
        RECT 96.980 192.430 97.300 193.630 ;
        RECT 94.420 191.230 96.660 191.630 ;
        RECT 97.620 190.870 101.820 209.910 ;
        RECT 103.420 208.930 105.660 209.330 ;
        RECT 102.140 206.930 102.460 208.130 ;
        RECT 102.780 207.330 105.020 207.730 ;
        RECT 105.980 206.930 106.300 208.130 ;
        RECT 103.420 205.730 105.660 206.130 ;
        RECT 103.420 201.430 105.660 201.830 ;
        RECT 102.140 199.430 102.460 200.630 ;
        RECT 102.780 199.830 105.020 200.230 ;
        RECT 105.980 199.430 106.300 200.630 ;
        RECT 103.420 198.230 105.660 198.630 ;
        RECT 103.420 194.430 105.660 194.830 ;
        RECT 102.140 192.430 102.460 193.630 ;
        RECT 102.780 192.830 105.020 193.230 ;
        RECT 105.980 192.430 106.300 193.630 ;
        RECT 103.420 191.230 105.660 191.630 ;
        RECT 106.620 190.870 107.580 209.910 ;
        RECT 10.460 189.910 107.580 190.870 ;
        RECT 109.020 195.030 109.660 210.950 ;
        RECT 110.840 208.990 112.280 210.190 ;
        RECT 111.920 205.390 112.280 208.990 ;
        RECT 113.000 208.990 114.440 210.190 ;
        RECT 113.000 205.390 113.360 208.990 ;
        RECT 114.080 205.390 114.440 208.990 ;
        RECT 115.160 208.990 116.600 210.190 ;
        RECT 115.160 205.390 115.520 208.990 ;
        RECT 111.920 195.790 113.360 198.190 ;
        RECT 114.080 195.790 115.520 198.190 ;
        RECT 117.780 195.030 119.020 210.950 ;
        RECT 109.020 192.950 119.020 195.030 ;
        RECT 43.520 189.890 56.020 189.910 ;
        RECT 61.520 189.890 74.020 189.910 ;
        RECT 13.020 187.890 35.520 188.890 ;
        RECT 13.020 172.030 13.660 187.890 ;
        RECT 14.840 185.990 16.280 187.190 ;
        RECT 15.920 182.390 16.280 185.990 ;
        RECT 17.000 185.990 18.440 187.190 ;
        RECT 17.000 182.390 17.360 185.990 ;
        RECT 18.080 182.390 18.440 185.990 ;
        RECT 19.160 185.990 20.600 187.190 ;
        RECT 19.160 182.390 19.520 185.990 ;
        RECT 20.240 182.390 20.600 185.990 ;
        RECT 21.320 185.990 22.760 187.190 ;
        RECT 21.320 182.390 21.680 185.990 ;
        RECT 22.400 182.390 22.760 185.990 ;
        RECT 23.480 185.990 24.920 187.190 ;
        RECT 23.480 182.390 23.840 185.990 ;
        RECT 24.560 182.390 24.920 185.990 ;
        RECT 25.640 185.990 27.080 187.190 ;
        RECT 25.640 182.390 26.000 185.990 ;
        RECT 26.720 182.390 27.080 185.990 ;
        RECT 27.800 185.990 29.240 187.190 ;
        RECT 27.800 182.390 28.160 185.990 ;
        RECT 28.880 182.390 29.240 185.990 ;
        RECT 29.960 185.990 31.400 187.190 ;
        RECT 29.960 182.390 30.320 185.990 ;
        RECT 31.040 182.390 31.400 185.990 ;
        RECT 32.120 185.990 33.560 187.190 ;
        RECT 32.120 182.390 32.480 185.990 ;
        RECT 15.920 172.790 17.360 175.190 ;
        RECT 18.080 172.790 19.520 175.190 ;
        RECT 20.240 172.790 21.680 175.190 ;
        RECT 22.400 172.790 23.840 175.190 ;
        RECT 24.560 172.790 26.000 175.190 ;
        RECT 26.720 172.790 28.160 175.190 ;
        RECT 28.880 172.790 30.320 175.190 ;
        RECT 31.040 172.790 32.480 175.190 ;
        RECT 34.740 172.870 35.520 187.890 ;
        RECT 82.740 188.390 104.940 188.510 ;
        RECT 109.020 188.390 109.660 192.950 ;
        RECT 110.840 190.990 112.280 192.190 ;
        RECT 82.740 187.950 109.660 188.390 ;
        RECT 37.460 186.910 53.180 187.870 ;
        RECT 37.460 174.870 38.420 186.910 ;
        RECT 39.380 185.930 41.620 186.330 ;
        RECT 38.740 183.930 39.060 185.130 ;
        RECT 40.020 184.330 42.260 184.730 ;
        RECT 42.580 183.930 42.900 185.130 ;
        RECT 39.380 182.730 41.620 183.130 ;
        RECT 39.380 178.430 41.620 178.830 ;
        RECT 38.740 176.430 39.060 177.630 ;
        RECT 40.020 176.830 42.260 177.230 ;
        RECT 42.580 176.430 42.900 177.630 ;
        RECT 39.380 175.230 41.620 175.630 ;
        RECT 43.220 174.870 47.420 186.910 ;
        RECT 48.380 185.430 50.620 185.830 ;
        RECT 47.740 183.430 48.060 184.630 ;
        RECT 49.020 183.830 51.260 184.230 ;
        RECT 51.580 183.430 51.900 184.630 ;
        RECT 48.380 182.230 50.620 182.630 ;
        RECT 48.380 178.430 50.620 178.830 ;
        RECT 47.740 176.430 48.060 177.630 ;
        RECT 49.020 176.830 51.260 177.230 ;
        RECT 51.580 176.430 51.900 177.630 ;
        RECT 48.380 175.230 50.620 175.630 ;
        RECT 52.220 174.870 53.180 186.910 ;
        RECT 37.460 173.910 53.180 174.870 ;
        RECT 64.860 186.910 80.580 187.870 ;
        RECT 64.860 174.870 65.820 186.910 ;
        RECT 67.420 185.430 69.660 185.830 ;
        RECT 66.140 183.430 66.460 184.630 ;
        RECT 66.780 183.830 69.020 184.230 ;
        RECT 69.980 183.430 70.300 184.630 ;
        RECT 67.420 182.230 69.660 182.630 ;
        RECT 67.420 178.430 69.660 178.830 ;
        RECT 66.140 176.430 66.460 177.630 ;
        RECT 66.780 176.830 69.020 177.230 ;
        RECT 69.980 176.430 70.300 177.630 ;
        RECT 67.420 175.230 69.660 175.630 ;
        RECT 70.620 174.870 74.820 186.910 ;
        RECT 76.420 185.930 78.660 186.330 ;
        RECT 75.140 183.930 75.460 185.130 ;
        RECT 75.780 184.330 78.020 184.730 ;
        RECT 78.980 183.930 79.300 185.130 ;
        RECT 76.420 182.730 78.660 183.130 ;
        RECT 76.420 178.430 78.660 178.830 ;
        RECT 75.140 176.430 75.460 177.630 ;
        RECT 75.780 176.830 78.020 177.230 ;
        RECT 78.980 176.430 79.300 177.630 ;
        RECT 76.420 175.230 78.660 175.630 ;
        RECT 79.620 174.870 80.580 186.910 ;
        RECT 64.860 173.910 80.580 174.870 ;
        RECT 34.740 172.390 80.580 172.870 ;
        RECT 82.740 172.390 83.300 187.950 ;
        RECT 84.480 185.990 85.920 187.190 ;
        RECT 85.560 182.390 85.920 185.990 ;
        RECT 86.640 185.990 88.080 187.190 ;
        RECT 86.640 182.390 87.000 185.990 ;
        RECT 87.720 182.390 88.080 185.990 ;
        RECT 88.800 185.990 90.240 187.190 ;
        RECT 88.800 182.390 89.160 185.990 ;
        RECT 89.880 182.390 90.240 185.990 ;
        RECT 90.960 185.990 92.400 187.190 ;
        RECT 90.960 182.390 91.320 185.990 ;
        RECT 92.040 182.390 92.400 185.990 ;
        RECT 93.120 185.990 94.560 187.190 ;
        RECT 93.120 182.390 93.480 185.990 ;
        RECT 94.200 182.390 94.560 185.990 ;
        RECT 95.280 185.990 96.720 187.190 ;
        RECT 95.280 182.390 95.640 185.990 ;
        RECT 96.360 182.390 96.720 185.990 ;
        RECT 97.440 185.990 98.880 187.190 ;
        RECT 97.440 182.390 97.800 185.990 ;
        RECT 98.520 182.390 98.880 185.990 ;
        RECT 99.600 185.990 101.040 187.190 ;
        RECT 99.600 182.390 99.960 185.990 ;
        RECT 100.680 182.390 101.040 185.990 ;
        RECT 101.760 185.990 103.200 187.190 ;
        RECT 101.760 182.390 102.120 185.990 ;
        RECT 104.380 177.030 109.660 187.950 ;
        RECT 111.920 187.390 112.280 190.990 ;
        RECT 113.000 190.990 114.440 192.190 ;
        RECT 113.000 187.390 113.360 190.990 ;
        RECT 114.080 187.390 114.440 190.990 ;
        RECT 115.160 190.990 116.600 192.190 ;
        RECT 115.160 187.390 115.520 190.990 ;
        RECT 111.920 177.790 113.360 180.190 ;
        RECT 114.080 177.790 115.520 180.190 ;
        RECT 117.780 177.030 119.020 192.950 ;
        RECT 85.560 172.790 87.000 175.190 ;
        RECT 87.720 172.790 89.160 175.190 ;
        RECT 89.880 172.790 91.320 175.190 ;
        RECT 92.040 172.790 93.480 175.190 ;
        RECT 94.200 172.790 95.640 175.190 ;
        RECT 96.360 172.790 97.800 175.190 ;
        RECT 98.520 172.790 99.960 175.190 ;
        RECT 100.680 172.790 102.120 175.190 ;
        RECT 104.380 174.950 119.020 177.030 ;
        RECT 34.740 172.030 83.300 172.390 ;
        RECT 104.380 172.030 109.660 174.950 ;
        RECT 110.840 172.990 112.280 174.190 ;
        RECT 13.020 171.910 109.660 172.030 ;
        RECT 13.020 169.950 38.420 171.910 ;
        RECT 39.380 170.430 41.620 170.830 ;
        RECT 13.020 154.030 13.660 169.950 ;
        RECT 32.360 169.190 33.560 169.950 ;
        RECT 14.840 167.990 16.280 169.190 ;
        RECT 15.920 164.390 16.280 167.990 ;
        RECT 17.000 167.990 18.440 169.190 ;
        RECT 17.000 164.390 17.360 167.990 ;
        RECT 18.080 164.390 18.440 167.990 ;
        RECT 19.160 167.990 20.600 169.190 ;
        RECT 19.160 164.390 19.520 167.990 ;
        RECT 20.240 164.390 20.600 167.990 ;
        RECT 21.320 167.990 22.760 169.190 ;
        RECT 21.320 164.390 21.680 167.990 ;
        RECT 22.400 164.390 22.760 167.990 ;
        RECT 23.480 167.990 24.920 169.190 ;
        RECT 23.480 164.390 23.840 167.990 ;
        RECT 24.560 164.390 24.920 167.990 ;
        RECT 25.640 167.990 27.080 169.190 ;
        RECT 25.640 164.390 26.000 167.990 ;
        RECT 26.720 164.390 27.080 167.990 ;
        RECT 27.800 167.990 29.240 169.190 ;
        RECT 27.800 164.390 28.160 167.990 ;
        RECT 28.880 164.390 29.240 167.990 ;
        RECT 29.960 167.990 31.400 169.190 ;
        RECT 29.960 164.390 30.320 167.990 ;
        RECT 31.040 164.390 31.400 167.990 ;
        RECT 32.120 167.990 33.560 169.190 ;
        RECT 32.120 164.390 32.480 167.990 ;
        RECT 34.740 161.890 38.420 169.950 ;
        RECT 38.740 168.430 39.060 169.630 ;
        RECT 40.020 168.830 42.260 169.230 ;
        RECT 42.580 168.430 42.900 169.630 ;
        RECT 39.380 167.230 41.620 167.630 ;
        RECT 39.380 165.430 41.620 165.830 ;
        RECT 38.740 163.430 39.060 164.630 ;
        RECT 40.020 163.830 42.260 164.230 ;
        RECT 42.580 163.430 42.900 164.630 ;
        RECT 39.380 162.230 41.620 162.630 ;
        RECT 43.220 161.890 47.420 171.910 ;
        RECT 48.380 170.430 50.620 170.830 ;
        RECT 47.740 168.430 48.060 169.630 ;
        RECT 49.020 168.830 51.260 169.230 ;
        RECT 51.580 168.430 51.900 169.630 ;
        RECT 48.380 167.230 50.620 167.630 ;
        RECT 48.380 165.430 50.620 165.830 ;
        RECT 47.740 163.430 48.060 164.630 ;
        RECT 49.020 163.830 51.260 164.230 ;
        RECT 51.580 163.430 51.900 164.630 ;
        RECT 48.380 162.230 50.620 162.630 ;
        RECT 52.220 161.890 65.820 171.910 ;
        RECT 67.420 170.430 69.660 170.830 ;
        RECT 66.140 168.430 66.460 169.630 ;
        RECT 66.780 168.830 69.020 169.230 ;
        RECT 69.980 168.430 70.300 169.630 ;
        RECT 67.420 167.230 69.660 167.630 ;
        RECT 67.420 165.430 69.660 165.830 ;
        RECT 66.140 163.430 66.460 164.630 ;
        RECT 66.780 163.830 69.020 164.230 ;
        RECT 69.980 163.430 70.300 164.630 ;
        RECT 67.420 162.230 69.660 162.630 ;
        RECT 34.740 161.870 65.820 161.890 ;
        RECT 70.620 161.870 74.820 171.910 ;
        RECT 76.420 170.430 78.660 170.830 ;
        RECT 79.620 169.950 109.660 171.910 ;
        RECT 75.140 168.430 75.460 169.630 ;
        RECT 75.780 168.830 78.020 169.230 ;
        RECT 78.980 168.430 79.300 169.630 ;
        RECT 76.420 167.230 78.660 167.630 ;
        RECT 76.420 165.430 78.660 165.830 ;
        RECT 75.140 163.430 75.460 164.630 ;
        RECT 75.780 163.830 78.020 164.230 ;
        RECT 78.980 163.430 79.300 164.630 ;
        RECT 76.420 162.230 78.660 162.630 ;
        RECT 79.620 161.870 83.300 169.950 ;
        RECT 84.480 169.190 85.680 169.950 ;
        RECT 84.480 167.990 85.920 169.190 ;
        RECT 85.560 164.390 85.920 167.990 ;
        RECT 86.640 167.990 88.080 169.190 ;
        RECT 86.640 164.390 87.000 167.990 ;
        RECT 87.720 164.390 88.080 167.990 ;
        RECT 88.800 167.990 90.240 169.190 ;
        RECT 88.800 164.390 89.160 167.990 ;
        RECT 89.880 164.390 90.240 167.990 ;
        RECT 90.960 167.990 92.400 169.190 ;
        RECT 90.960 164.390 91.320 167.990 ;
        RECT 92.040 164.390 92.400 167.990 ;
        RECT 93.120 167.990 94.560 169.190 ;
        RECT 93.120 164.390 93.480 167.990 ;
        RECT 94.200 164.390 94.560 167.990 ;
        RECT 95.280 167.990 96.720 169.190 ;
        RECT 95.280 164.390 95.640 167.990 ;
        RECT 96.360 164.390 96.720 167.990 ;
        RECT 97.440 167.990 98.880 169.190 ;
        RECT 97.440 164.390 97.800 167.990 ;
        RECT 98.520 164.390 98.880 167.990 ;
        RECT 99.600 167.990 101.040 169.190 ;
        RECT 99.600 164.390 99.960 167.990 ;
        RECT 100.680 164.390 101.040 167.990 ;
        RECT 101.760 167.990 103.200 169.190 ;
        RECT 101.760 164.390 102.120 167.990 ;
        RECT 34.740 160.910 83.300 161.870 ;
        RECT 34.740 160.390 65.520 160.910 ;
        RECT 15.920 154.790 17.360 157.190 ;
        RECT 18.080 154.790 19.520 157.190 ;
        RECT 20.240 154.790 21.680 157.190 ;
        RECT 22.400 154.790 23.840 157.190 ;
        RECT 24.560 154.790 26.000 157.190 ;
        RECT 26.720 154.790 28.160 157.190 ;
        RECT 28.880 154.790 30.320 157.190 ;
        RECT 31.040 154.790 32.480 157.190 ;
        RECT 34.740 156.785 61.020 160.390 ;
        RECT 63.120 157.770 64.020 158.990 ;
        RECT 65.970 158.240 70.320 158.540 ;
        RECT 64.920 157.840 65.820 158.140 ;
        RECT 71.220 157.840 72.120 158.140 ;
        RECT 61.940 156.810 64.020 157.770 ;
        RECT 66.780 157.740 67.620 157.760 ;
        RECT 69.480 157.740 70.320 157.760 ;
        RECT 66.720 157.440 67.620 157.740 ;
        RECT 69.420 157.440 70.320 157.740 ;
        RECT 70.620 157.540 71.520 157.840 ;
        RECT 73.020 157.730 73.920 158.990 ;
        RECT 64.920 157.040 65.820 157.340 ;
        RECT 70.620 157.240 70.920 157.540 ;
        RECT 70.020 156.940 70.920 157.240 ;
        RECT 71.220 157.040 72.570 157.340 ;
        RECT 34.740 154.030 39.325 156.785 ;
        RECT 13.020 152.695 39.325 154.030 ;
        RECT 39.635 153.005 43.105 156.475 ;
        RECT 43.415 152.695 47.325 156.785 ;
        RECT 47.635 153.005 51.105 156.475 ;
        RECT 51.415 152.695 55.325 156.785 ;
        RECT 55.635 153.005 59.105 156.475 ;
        RECT 59.415 154.390 61.020 156.785 ;
        RECT 63.120 156.190 64.020 156.810 ;
        RECT 66.720 156.640 70.320 156.940 ;
        RECT 73.020 156.850 75.160 157.730 ;
        RECT 73.020 156.190 73.920 156.850 ;
        RECT 74.280 155.450 75.160 156.850 ;
        RECT 59.415 153.890 63.020 154.390 ;
        RECT 59.415 152.695 63.220 153.890 ;
        RECT 67.870 153.440 68.170 154.040 ;
        RECT 80.520 154.030 83.300 160.910 ;
        RECT 104.380 159.030 109.660 169.950 ;
        RECT 111.920 169.390 112.280 172.990 ;
        RECT 113.000 172.990 114.440 174.190 ;
        RECT 113.000 169.390 113.360 172.990 ;
        RECT 114.080 169.390 114.440 172.990 ;
        RECT 115.160 172.990 116.600 174.190 ;
        RECT 115.160 169.390 115.520 172.990 ;
        RECT 111.920 159.790 113.360 162.190 ;
        RECT 114.080 159.790 115.520 162.190 ;
        RECT 117.780 159.030 119.020 174.950 ;
        RECT 85.560 154.790 87.000 157.190 ;
        RECT 87.720 154.790 89.160 157.190 ;
        RECT 89.880 154.790 91.320 157.190 ;
        RECT 92.040 154.790 93.480 157.190 ;
        RECT 94.200 154.790 95.640 157.190 ;
        RECT 96.360 154.790 97.800 157.190 ;
        RECT 98.520 154.790 99.960 157.190 ;
        RECT 100.680 154.790 102.120 157.190 ;
        RECT 104.380 156.950 119.020 159.030 ;
        RECT 104.380 156.190 109.660 156.950 ;
        RECT 104.380 154.990 112.280 156.190 ;
        RECT 104.380 154.030 109.660 154.990 ;
        RECT 68.620 153.440 69.460 153.460 ;
        RECT 65.920 153.140 69.520 153.440 ;
        RECT 64.120 152.740 65.620 153.040 ;
        RECT 70.420 152.740 71.320 153.040 ;
        RECT 13.020 151.890 63.220 152.695 ;
        RECT 13.020 136.030 13.660 151.890 ;
        RECT 14.840 149.990 16.280 151.190 ;
        RECT 15.920 146.390 16.280 149.990 ;
        RECT 17.000 149.990 18.440 151.190 ;
        RECT 17.000 146.390 17.360 149.990 ;
        RECT 18.080 146.390 18.440 149.990 ;
        RECT 19.160 149.990 20.600 151.190 ;
        RECT 19.160 146.390 19.520 149.990 ;
        RECT 20.240 146.390 20.600 149.990 ;
        RECT 21.320 149.990 22.760 151.190 ;
        RECT 21.320 146.390 21.680 149.990 ;
        RECT 22.400 146.390 22.760 149.990 ;
        RECT 23.480 149.990 24.920 151.190 ;
        RECT 23.480 146.390 23.840 149.990 ;
        RECT 24.560 146.390 24.920 149.990 ;
        RECT 25.640 149.990 27.080 151.190 ;
        RECT 25.640 146.390 26.000 149.990 ;
        RECT 26.720 146.390 27.080 149.990 ;
        RECT 27.800 149.990 29.240 151.190 ;
        RECT 27.800 146.390 28.160 149.990 ;
        RECT 28.880 146.390 29.240 149.990 ;
        RECT 29.960 149.990 31.400 151.190 ;
        RECT 29.960 146.390 30.320 149.990 ;
        RECT 31.040 146.390 31.400 149.990 ;
        RECT 32.120 149.990 33.560 151.190 ;
        RECT 32.120 146.390 32.480 149.990 ;
        RECT 34.740 148.785 63.220 151.890 ;
        RECT 65.320 151.840 65.620 152.740 ;
        RECT 65.920 152.640 66.760 152.660 ;
        RECT 68.620 152.640 69.460 152.660 ;
        RECT 65.920 152.340 66.820 152.640 ;
        RECT 68.620 152.340 69.520 152.640 ;
        RECT 65.920 151.840 66.760 151.860 ;
        RECT 65.320 151.540 69.520 151.840 ;
        RECT 64.120 151.440 64.960 151.460 ;
        RECT 64.120 151.140 65.020 151.440 ;
        RECT 69.820 151.140 71.320 151.440 ;
        RECT 65.920 150.740 69.520 151.040 ;
        RECT 64.120 150.340 65.020 150.640 ;
        RECT 65.920 149.940 66.820 150.240 ;
        RECT 64.120 149.840 64.960 149.860 ;
        RECT 64.120 149.540 65.020 149.840 ;
        RECT 65.920 149.440 66.760 149.460 ;
        RECT 68.020 149.440 68.320 150.740 ;
        RECT 68.620 150.240 69.460 150.260 ;
        RECT 68.620 149.940 69.520 150.240 ;
        RECT 65.920 149.140 66.820 149.440 ;
        RECT 68.020 149.140 69.520 149.440 ;
        RECT 34.740 144.695 39.325 148.785 ;
        RECT 39.635 145.005 43.105 148.475 ;
        RECT 43.415 144.695 47.325 148.785 ;
        RECT 47.635 145.005 51.105 148.475 ;
        RECT 51.415 144.695 55.325 148.785 ;
        RECT 55.635 145.005 59.105 148.475 ;
        RECT 59.415 144.695 63.220 148.785 ;
        RECT 65.920 148.640 66.760 148.660 ;
        RECT 65.920 148.340 69.520 148.640 ;
        RECT 64.120 147.940 65.020 148.240 ;
        RECT 64.720 147.640 65.620 147.940 ;
        RECT 64.120 147.140 65.020 147.440 ;
        RECT 64.120 145.840 64.960 145.860 ;
        RECT 64.120 145.540 65.020 145.840 ;
        RECT 34.740 140.785 63.220 144.695 ;
        RECT 65.320 144.240 65.620 147.640 ;
        RECT 65.920 147.540 66.820 147.840 ;
        RECT 68.620 147.540 69.520 147.840 ;
        RECT 65.920 147.040 66.760 147.060 ;
        RECT 68.620 147.040 69.460 147.060 ;
        RECT 65.920 146.740 66.820 147.040 ;
        RECT 68.620 146.740 69.520 147.040 ;
        RECT 68.620 146.240 69.460 146.260 ;
        RECT 65.920 145.940 69.520 146.240 ;
        RECT 65.920 145.440 66.760 145.460 ;
        RECT 68.620 145.440 69.460 145.460 ;
        RECT 65.920 145.140 66.820 145.440 ;
        RECT 68.620 145.140 69.520 145.440 ;
        RECT 65.920 144.640 66.760 144.660 ;
        RECT 65.920 144.340 69.520 144.640 ;
        RECT 64.120 143.940 65.620 144.240 ;
        RECT 64.120 143.140 65.020 143.440 ;
        RECT 64.120 141.840 64.960 141.860 ;
        RECT 64.120 141.540 65.020 141.840 ;
        RECT 15.920 136.790 17.360 139.190 ;
        RECT 18.080 136.790 19.520 139.190 ;
        RECT 20.240 136.790 21.680 139.190 ;
        RECT 22.400 136.790 23.840 139.190 ;
        RECT 24.560 136.790 26.000 139.190 ;
        RECT 26.720 136.790 28.160 139.190 ;
        RECT 28.880 136.790 30.320 139.190 ;
        RECT 31.040 136.790 32.480 139.190 ;
        RECT 34.740 136.695 39.325 140.785 ;
        RECT 39.635 137.005 43.105 140.475 ;
        RECT 43.415 136.695 47.325 140.785 ;
        RECT 47.635 137.005 51.105 140.475 ;
        RECT 51.415 136.695 55.325 140.785 ;
        RECT 55.635 137.005 59.105 140.475 ;
        RECT 59.415 136.695 63.220 140.785 ;
        RECT 64.120 140.740 65.020 141.040 ;
        RECT 65.320 139.840 65.620 143.940 ;
        RECT 65.920 143.540 66.820 143.840 ;
        RECT 65.920 143.040 66.760 143.060 ;
        RECT 65.920 142.740 66.820 143.040 ;
        RECT 67.120 142.240 67.420 144.340 ;
        RECT 68.620 143.540 69.520 143.840 ;
        RECT 68.620 143.040 69.460 143.060 ;
        RECT 68.620 142.740 69.520 143.040 ;
        RECT 65.920 141.940 69.520 142.240 ;
        RECT 69.820 141.840 70.120 151.140 ;
        RECT 70.420 150.640 71.260 150.660 ;
        RECT 70.420 150.340 71.320 150.640 ;
        RECT 70.420 149.540 71.320 149.840 ;
        RECT 70.420 148.240 71.260 148.260 ;
        RECT 70.420 147.940 71.320 148.240 ;
        RECT 70.420 147.440 71.260 147.460 ;
        RECT 70.420 147.140 71.320 147.440 ;
        RECT 70.420 145.540 71.320 145.840 ;
        RECT 70.420 144.240 71.260 144.260 ;
        RECT 70.420 143.940 71.320 144.240 ;
        RECT 70.420 143.440 71.260 143.460 ;
        RECT 70.420 143.140 71.320 143.440 ;
        RECT 69.820 141.540 71.320 141.840 ;
        RECT 65.920 141.140 66.820 141.440 ;
        RECT 68.620 141.140 69.520 141.440 ;
        RECT 65.920 140.640 66.760 140.660 ;
        RECT 68.620 140.640 69.460 140.660 ;
        RECT 65.920 140.340 66.820 140.640 ;
        RECT 68.620 140.340 69.520 140.640 ;
        RECT 69.820 139.840 70.120 141.540 ;
        RECT 70.420 140.740 71.320 141.040 ;
        RECT 70.870 140.240 71.170 140.740 ;
        RECT 65.320 139.540 70.120 139.840 ;
        RECT 64.120 139.140 65.020 139.440 ;
        RECT 70.420 139.140 71.320 139.440 ;
        RECT 65.920 139.040 66.760 139.060 ;
        RECT 68.620 139.040 69.460 139.060 ;
        RECT 65.920 138.740 66.820 139.040 ;
        RECT 68.620 138.740 69.520 139.040 ;
        RECT 69.820 138.840 70.720 139.140 ;
        RECT 65.920 138.240 66.760 138.260 ;
        RECT 68.620 138.240 69.460 138.260 ;
        RECT 65.920 137.940 67.420 138.240 ;
        RECT 68.620 137.940 69.520 138.240 ;
        RECT 64.120 137.840 64.960 137.860 ;
        RECT 64.120 137.540 65.020 137.840 ;
        RECT 67.120 137.440 67.420 137.940 ;
        RECT 68.620 137.440 69.460 137.460 ;
        RECT 69.820 137.440 70.120 138.840 ;
        RECT 70.420 137.540 71.320 137.840 ;
        RECT 65.920 137.140 66.820 137.440 ;
        RECT 67.120 137.140 70.120 137.440 ;
        RECT 63.870 136.740 65.020 137.040 ;
        RECT 70.420 136.740 71.320 137.040 ;
        RECT 34.740 136.030 63.220 136.695 ;
        RECT 65.920 136.640 66.760 136.660 ;
        RECT 68.620 136.640 69.460 136.660 ;
        RECT 65.920 136.340 66.820 136.640 ;
        RECT 68.620 136.340 69.520 136.640 ;
        RECT 13.020 135.440 63.220 136.030 ;
        RECT 65.920 135.840 66.760 135.860 ;
        RECT 68.620 135.840 69.460 135.860 ;
        RECT 65.320 135.540 66.820 135.840 ;
        RECT 68.620 135.540 70.120 135.840 ;
        RECT 65.320 135.440 65.620 135.540 ;
        RECT 13.020 135.140 65.620 135.440 ;
        RECT 13.020 134.290 63.220 135.140 ;
        RECT 65.320 135.040 65.620 135.140 ;
        RECT 69.820 135.440 70.120 135.540 ;
        RECT 72.220 135.440 73.120 153.890 ;
        RECT 80.520 153.390 109.660 154.030 ;
        RECT 69.820 135.140 73.120 135.440 ;
        RECT 65.920 135.040 66.760 135.060 ;
        RECT 68.620 135.040 69.460 135.060 ;
        RECT 69.820 135.040 70.120 135.140 ;
        RECT 65.320 134.740 66.820 135.040 ;
        RECT 68.620 134.740 70.120 135.040 ;
        RECT 13.020 133.890 63.020 134.290 ;
        RECT 13.020 118.030 13.660 133.890 ;
        RECT 14.840 131.990 16.280 133.190 ;
        RECT 15.920 128.390 16.280 131.990 ;
        RECT 17.000 131.990 18.440 133.190 ;
        RECT 17.000 128.390 17.360 131.990 ;
        RECT 18.080 128.390 18.440 131.990 ;
        RECT 19.160 131.990 20.600 133.190 ;
        RECT 19.160 128.390 19.520 131.990 ;
        RECT 20.240 128.390 20.600 131.990 ;
        RECT 21.320 131.990 22.760 133.190 ;
        RECT 21.320 128.390 21.680 131.990 ;
        RECT 22.400 128.390 22.760 131.990 ;
        RECT 23.480 131.990 24.920 133.190 ;
        RECT 23.480 128.390 23.840 131.990 ;
        RECT 24.560 128.390 24.920 131.990 ;
        RECT 25.640 131.990 27.080 133.190 ;
        RECT 25.640 128.390 26.000 131.990 ;
        RECT 26.720 128.390 27.080 131.990 ;
        RECT 27.800 131.990 29.240 133.190 ;
        RECT 27.800 128.390 28.160 131.990 ;
        RECT 28.880 128.390 29.240 131.990 ;
        RECT 29.960 131.990 31.400 133.190 ;
        RECT 29.960 128.390 30.320 131.990 ;
        RECT 31.040 128.390 31.400 131.990 ;
        RECT 32.120 131.990 33.560 133.190 ;
        RECT 32.120 128.390 32.480 131.990 ;
        RECT 15.920 118.790 17.360 121.190 ;
        RECT 18.080 118.790 19.520 121.190 ;
        RECT 20.240 118.790 21.680 121.190 ;
        RECT 22.400 118.790 23.840 121.190 ;
        RECT 24.560 118.790 26.000 121.190 ;
        RECT 26.720 118.790 28.160 121.190 ;
        RECT 28.880 118.790 30.320 121.190 ;
        RECT 31.040 118.790 32.480 121.190 ;
        RECT 34.740 118.030 37.660 133.890 ;
        RECT 38.840 131.990 40.280 133.190 ;
        RECT 39.920 128.390 40.280 131.990 ;
        RECT 41.000 131.990 42.440 133.190 ;
        RECT 41.000 128.390 41.360 131.990 ;
        RECT 42.080 128.390 42.440 131.990 ;
        RECT 43.160 131.990 44.600 133.190 ;
        RECT 43.160 128.390 43.520 131.990 ;
        RECT 44.240 128.390 44.600 131.990 ;
        RECT 45.320 131.990 46.760 133.190 ;
        RECT 45.320 128.390 45.680 131.990 ;
        RECT 46.400 128.390 46.760 131.990 ;
        RECT 47.480 131.990 48.920 133.190 ;
        RECT 47.480 128.390 47.840 131.990 ;
        RECT 48.560 128.390 48.920 131.990 ;
        RECT 49.640 131.990 51.080 133.190 ;
        RECT 49.640 128.390 50.000 131.990 ;
        RECT 50.720 128.390 51.080 131.990 ;
        RECT 51.800 131.990 53.240 133.190 ;
        RECT 51.800 128.390 52.160 131.990 ;
        RECT 52.880 128.390 53.240 131.990 ;
        RECT 53.960 131.990 55.400 133.190 ;
        RECT 53.960 128.390 54.320 131.990 ;
        RECT 55.040 128.390 55.400 131.990 ;
        RECT 56.120 131.990 57.560 133.190 ;
        RECT 56.120 128.390 56.480 131.990 ;
        RECT 58.740 124.370 60.920 133.890 ;
        RECT 69.670 133.840 69.970 134.740 ;
        RECT 72.220 134.290 73.120 135.140 ;
        RECT 77.020 141.030 109.660 153.390 ;
        RECT 111.920 151.390 112.280 154.990 ;
        RECT 113.000 154.990 114.440 156.190 ;
        RECT 113.000 151.390 113.360 154.990 ;
        RECT 114.080 151.390 114.440 154.990 ;
        RECT 115.160 154.990 116.600 156.190 ;
        RECT 115.160 151.390 115.520 154.990 ;
        RECT 111.920 141.790 113.360 144.190 ;
        RECT 114.080 141.790 115.520 144.190 ;
        RECT 117.780 141.030 119.020 156.950 ;
        RECT 77.020 139.890 119.020 141.030 ;
        RECT 77.020 136.390 105.020 139.890 ;
        RECT 65.080 132.890 66.040 133.530 ;
        RECT 77.020 132.890 85.520 136.390 ;
        RECT 61.880 131.930 63.480 132.330 ;
        RECT 61.240 130.730 61.560 131.930 ;
        RECT 62.520 131.130 64.120 131.530 ;
        RECT 64.440 130.730 64.760 131.930 ;
        RECT 61.880 130.330 63.480 130.730 ;
        RECT 61.880 127.130 63.480 127.530 ;
        RECT 61.240 125.930 61.560 127.130 ;
        RECT 62.520 126.330 64.120 126.730 ;
        RECT 64.440 125.930 64.760 127.130 ;
        RECT 61.880 125.530 63.480 125.930 ;
        RECT 65.080 124.370 85.520 132.890 ;
        RECT 58.740 121.890 85.520 124.370 ;
        RECT 39.920 118.790 41.360 121.190 ;
        RECT 42.080 118.790 43.520 121.190 ;
        RECT 44.240 118.790 45.680 121.190 ;
        RECT 46.400 118.790 47.840 121.190 ;
        RECT 48.560 118.790 50.000 121.190 ;
        RECT 50.720 118.790 52.160 121.190 ;
        RECT 52.880 118.790 54.320 121.190 ;
        RECT 55.040 118.790 56.480 121.190 ;
        RECT 58.740 118.030 59.520 121.890 ;
        RECT 13.020 117.390 59.520 118.030 ;
        RECT 74.180 96.170 75.140 101.600 ;
        RECT 76.100 99.530 78.340 99.930 ;
        RECT 75.460 97.530 75.780 98.730 ;
        RECT 76.740 97.930 78.980 98.330 ;
        RECT 79.300 97.530 79.620 98.730 ;
        RECT 76.100 96.330 78.340 96.730 ;
        RECT 79.940 96.170 80.900 101.600 ;
        RECT 91.230 101.550 121.060 101.710 ;
        RECT 74.160 95.930 75.140 96.170 ;
        RECT 79.920 95.930 80.900 96.170 ;
        RECT 90.560 101.150 121.060 101.550 ;
        RECT 90.560 100.990 99.800 101.150 ;
        RECT 63.020 90.280 63.980 94.410 ;
        RECT 64.940 93.610 67.180 94.010 ;
        RECT 64.300 91.610 64.620 92.810 ;
        RECT 65.580 92.010 67.820 92.410 ;
        RECT 68.140 91.610 68.460 92.810 ;
        RECT 64.940 90.410 67.180 90.810 ;
        RECT 68.780 90.280 69.740 94.410 ;
        RECT 74.160 92.180 75.120 95.930 ;
        RECT 76.080 95.370 78.320 95.770 ;
        RECT 75.440 93.370 75.760 94.570 ;
        RECT 76.720 93.770 78.960 94.170 ;
        RECT 79.280 93.370 79.600 94.570 ;
        RECT 74.160 91.770 75.160 92.180 ;
        RECT 76.080 92.170 78.320 92.570 ;
        RECT 79.920 92.180 80.880 95.930 ;
        RECT 63.010 90.010 63.980 90.280 ;
        RECT 68.770 90.010 69.740 90.280 ;
        RECT 63.010 86.280 63.970 90.010 ;
        RECT 64.930 89.480 67.170 89.880 ;
        RECT 64.290 87.480 64.610 88.680 ;
        RECT 65.570 87.880 67.810 88.280 ;
        RECT 68.130 87.480 68.450 88.680 ;
        RECT 64.930 86.280 67.170 86.680 ;
        RECT 68.770 86.280 69.730 90.010 ;
        RECT 74.200 88.020 75.160 91.770 ;
        RECT 76.120 91.380 78.360 91.780 ;
        RECT 79.920 91.770 80.920 92.180 ;
        RECT 75.480 89.380 75.800 90.580 ;
        RECT 76.760 89.780 79.000 90.180 ;
        RECT 79.320 89.380 79.640 90.580 ;
        RECT 76.120 88.180 78.360 88.580 ;
        RECT 79.960 88.020 80.920 91.770 ;
        RECT 74.160 87.780 75.160 88.020 ;
        RECT 79.920 87.780 80.920 88.020 ;
        RECT 63.010 85.880 64.000 86.280 ;
        RECT 68.770 85.880 69.760 86.280 ;
        RECT 63.040 82.150 64.000 85.880 ;
        RECT 64.960 85.480 67.200 85.880 ;
        RECT 64.320 83.480 64.640 84.680 ;
        RECT 65.600 83.880 67.840 84.280 ;
        RECT 68.160 83.480 68.480 84.680 ;
        RECT 64.960 82.280 67.200 82.680 ;
        RECT 68.800 82.150 69.760 85.880 ;
        RECT 74.160 84.020 75.120 87.780 ;
        RECT 76.080 87.220 78.320 87.620 ;
        RECT 75.440 85.220 75.760 86.420 ;
        RECT 76.720 85.620 78.960 86.020 ;
        RECT 79.280 85.220 79.600 86.420 ;
        RECT 76.080 84.020 78.320 84.420 ;
        RECT 79.920 84.020 80.880 87.780 ;
        RECT 90.560 85.070 91.120 100.990 ;
        RECT 91.680 99.030 93.740 100.230 ;
        RECT 93.380 95.430 93.740 99.030 ;
        RECT 94.460 99.030 95.900 100.230 ;
        RECT 94.460 95.430 94.820 99.030 ;
        RECT 95.540 95.430 95.900 99.030 ;
        RECT 96.620 99.030 98.590 100.230 ;
        RECT 96.620 95.430 96.980 99.030 ;
        RECT 93.380 85.830 94.820 88.230 ;
        RECT 95.540 85.830 96.980 88.230 ;
        RECT 99.240 85.070 99.800 100.990 ;
        RECT 90.560 84.720 99.800 85.070 ;
        RECT 101.230 101.070 110.470 101.150 ;
        RECT 101.230 85.150 101.790 101.070 ;
        RECT 102.330 99.110 104.410 100.310 ;
        RECT 104.050 95.510 104.410 99.110 ;
        RECT 105.130 99.110 106.570 100.310 ;
        RECT 105.130 95.510 105.490 99.110 ;
        RECT 106.210 95.510 106.570 99.110 ;
        RECT 107.290 99.110 109.370 100.310 ;
        RECT 107.290 95.510 107.650 99.110 ;
        RECT 104.050 85.910 105.490 88.310 ;
        RECT 106.210 85.910 107.650 88.310 ;
        RECT 109.910 85.150 110.470 101.070 ;
        RECT 101.230 84.720 110.470 85.150 ;
        RECT 111.820 85.230 112.380 101.150 ;
        RECT 118.060 100.390 119.260 101.150 ;
        RECT 112.950 99.190 115.000 100.390 ;
        RECT 114.640 95.590 115.000 99.190 ;
        RECT 115.720 99.190 117.160 100.390 ;
        RECT 115.720 95.590 116.080 99.190 ;
        RECT 116.800 95.590 117.160 99.190 ;
        RECT 117.880 99.190 119.990 100.390 ;
        RECT 117.880 95.590 118.240 99.190 ;
        RECT 114.640 85.990 116.080 88.390 ;
        RECT 116.800 85.990 118.240 88.390 ;
        RECT 120.500 85.230 121.060 101.150 ;
        RECT 111.820 84.720 121.060 85.230 ;
        RECT 90.560 84.510 159.340 84.720 ;
        RECT 74.160 83.620 75.140 84.020 ;
        RECT 79.920 83.620 80.900 84.020 ;
        RECT 63.030 81.880 64.000 82.150 ;
        RECT 68.790 81.880 69.760 82.150 ;
        RECT 63.030 78.160 63.990 81.880 ;
        RECT 64.950 81.350 67.190 81.750 ;
        RECT 64.310 79.350 64.630 80.550 ;
        RECT 65.590 79.750 67.830 80.150 ;
        RECT 68.150 79.350 68.470 80.550 ;
        RECT 63.030 77.750 64.000 78.160 ;
        RECT 64.950 78.150 67.190 78.550 ;
        RECT 68.790 78.160 69.750 81.880 ;
        RECT 74.180 79.860 75.140 83.620 ;
        RECT 76.100 83.220 78.340 83.620 ;
        RECT 75.460 81.220 75.780 82.420 ;
        RECT 76.740 81.620 78.980 82.020 ;
        RECT 79.300 81.220 79.620 82.420 ;
        RECT 76.100 80.020 78.340 80.420 ;
        RECT 79.940 79.860 80.900 83.620 ;
        RECT 74.160 79.620 75.140 79.860 ;
        RECT 79.920 79.620 80.900 79.860 ;
        RECT 63.040 74.030 64.000 77.750 ;
        RECT 64.960 77.360 67.200 77.760 ;
        RECT 68.790 77.750 69.760 78.160 ;
        RECT 64.320 75.360 64.640 76.560 ;
        RECT 65.600 75.760 67.840 76.160 ;
        RECT 68.160 75.360 68.480 76.560 ;
        RECT 64.960 74.160 67.200 74.560 ;
        RECT 68.800 74.030 69.760 77.750 ;
        RECT 74.160 75.730 75.120 79.620 ;
        RECT 76.080 79.060 78.320 79.460 ;
        RECT 75.440 77.060 75.760 78.260 ;
        RECT 76.720 77.460 78.960 77.860 ;
        RECT 79.280 77.060 79.600 78.260 ;
        RECT 76.080 75.860 78.320 76.260 ;
        RECT 79.920 75.730 80.880 79.620 ;
        RECT 90.690 76.620 159.340 84.510 ;
        RECT 92.580 76.150 159.340 76.620 ;
        RECT 74.160 75.460 75.140 75.730 ;
        RECT 79.920 75.460 80.900 75.730 ;
        RECT 63.030 73.760 64.000 74.030 ;
        RECT 68.790 73.760 69.760 74.030 ;
        RECT 35.700 72.870 36.660 72.890 ;
        RECT 4.650 72.670 26.850 72.780 ;
        RECT 33.780 72.770 40.530 72.870 ;
        RECT 0.470 72.220 26.850 72.670 ;
        RECT 0.470 56.300 5.300 72.220 ;
        RECT 6.390 70.260 7.830 71.460 ;
        RECT 7.470 66.660 7.830 70.260 ;
        RECT 8.550 70.260 9.990 71.460 ;
        RECT 8.550 66.660 8.910 70.260 ;
        RECT 9.630 66.660 9.990 70.260 ;
        RECT 10.710 70.260 12.150 71.460 ;
        RECT 10.710 66.660 11.070 70.260 ;
        RECT 11.790 66.660 12.150 70.260 ;
        RECT 12.870 70.260 14.310 71.460 ;
        RECT 12.870 66.660 13.230 70.260 ;
        RECT 13.950 66.660 14.310 70.260 ;
        RECT 15.030 70.260 16.470 71.460 ;
        RECT 15.030 66.660 15.390 70.260 ;
        RECT 16.110 66.660 16.470 70.260 ;
        RECT 17.190 70.260 18.630 71.460 ;
        RECT 17.190 66.660 17.550 70.260 ;
        RECT 18.270 66.660 18.630 70.260 ;
        RECT 19.350 70.260 20.790 71.460 ;
        RECT 19.350 66.660 19.710 70.260 ;
        RECT 20.430 66.660 20.790 70.260 ;
        RECT 21.510 70.260 22.950 71.460 ;
        RECT 21.510 66.660 21.870 70.260 ;
        RECT 22.590 66.660 22.950 70.260 ;
        RECT 23.670 70.260 25.110 71.460 ;
        RECT 23.670 66.660 24.030 70.260 ;
        RECT 7.470 57.060 8.910 59.460 ;
        RECT 9.630 57.060 11.070 59.460 ;
        RECT 11.790 57.060 13.230 59.460 ;
        RECT 13.950 57.060 15.390 59.460 ;
        RECT 16.110 57.060 17.550 59.460 ;
        RECT 18.270 57.060 19.710 59.460 ;
        RECT 20.430 57.060 21.870 59.460 ;
        RECT 22.590 57.060 24.030 59.460 ;
        RECT 26.290 56.300 26.850 72.220 ;
        RECT 33.770 71.910 40.530 72.770 ;
        RECT 33.770 71.810 40.500 71.910 ;
        RECT 33.780 68.770 34.740 71.810 ;
        RECT 35.700 68.910 36.660 71.810 ;
        RECT 39.540 68.770 40.500 71.810 ;
        RECT 63.030 70.020 63.990 73.760 ;
        RECT 64.950 73.230 67.190 73.630 ;
        RECT 64.310 71.230 64.630 72.430 ;
        RECT 65.590 71.630 67.830 72.030 ;
        RECT 68.150 71.230 68.470 72.430 ;
        RECT 64.950 70.030 67.190 70.430 ;
        RECT 68.790 70.020 69.750 73.760 ;
        RECT 74.180 71.570 75.140 75.460 ;
        RECT 76.100 74.930 78.340 75.330 ;
        RECT 75.460 72.930 75.780 74.130 ;
        RECT 76.740 73.330 78.980 73.730 ;
        RECT 79.300 72.930 79.620 74.130 ;
        RECT 76.100 71.730 78.340 72.130 ;
        RECT 79.940 71.570 80.900 75.460 ;
        RECT 74.180 71.330 75.150 71.570 ;
        RECT 79.940 71.330 80.910 71.570 ;
        RECT 63.030 69.630 64.020 70.020 ;
        RECT 68.790 69.630 69.780 70.020 ;
        RECT 33.770 67.620 34.740 68.770 ;
        RECT 35.690 67.970 37.930 68.370 ;
        RECT 33.770 64.860 34.730 67.620 ;
        RECT 39.530 67.390 40.500 68.770 ;
        RECT 35.050 65.970 35.370 67.170 ;
        RECT 36.330 66.370 38.570 66.770 ;
        RECT 38.890 65.970 39.210 67.170 ;
        RECT 33.770 64.370 34.760 64.860 ;
        RECT 35.690 64.770 37.930 65.170 ;
        RECT 39.530 65.140 40.490 67.390 ;
        RECT 63.060 65.890 64.020 69.630 ;
        RECT 64.980 69.220 67.220 69.620 ;
        RECT 64.340 67.220 64.660 68.420 ;
        RECT 65.620 67.620 67.860 68.020 ;
        RECT 68.180 67.220 68.500 68.420 ;
        RECT 64.980 66.020 67.220 66.420 ;
        RECT 68.820 65.890 69.780 69.630 ;
        RECT 74.190 67.440 75.150 71.330 ;
        RECT 76.110 70.770 78.350 71.170 ;
        RECT 75.470 68.770 75.790 69.970 ;
        RECT 76.750 69.170 78.990 69.570 ;
        RECT 79.310 68.770 79.630 69.970 ;
        RECT 76.110 67.570 78.350 67.970 ;
        RECT 79.950 67.440 80.910 71.330 ;
        RECT 63.050 65.620 64.020 65.890 ;
        RECT 68.810 65.620 69.780 65.890 ;
        RECT 74.170 67.170 75.150 67.440 ;
        RECT 79.930 67.170 80.910 67.440 ;
        RECT 39.530 64.370 40.520 65.140 ;
        RECT 33.800 63.750 34.760 64.370 ;
        RECT 39.560 63.750 40.520 64.370 ;
        RECT 33.790 62.020 34.760 63.750 ;
        RECT 35.710 62.950 37.950 63.350 ;
        RECT 33.790 59.350 34.750 62.020 ;
        RECT 35.070 60.950 35.390 62.150 ;
        RECT 36.350 61.350 38.590 61.750 ;
        RECT 38.910 60.950 39.230 62.150 ;
        RECT 39.550 62.040 40.520 63.750 ;
        RECT 35.710 59.750 37.950 60.150 ;
        RECT 39.550 59.350 40.510 62.040 ;
        RECT 63.050 61.900 64.010 65.620 ;
        RECT 64.970 65.090 67.210 65.490 ;
        RECT 64.330 63.090 64.650 64.290 ;
        RECT 65.610 63.490 67.850 63.890 ;
        RECT 68.170 63.090 68.490 64.290 ;
        RECT 63.050 61.490 64.020 61.900 ;
        RECT 64.970 61.890 67.210 62.290 ;
        RECT 68.810 61.900 69.770 65.620 ;
        RECT 74.170 63.280 75.130 67.170 ;
        RECT 76.090 66.640 78.330 67.040 ;
        RECT 75.450 64.640 75.770 65.840 ;
        RECT 76.730 65.040 78.970 65.440 ;
        RECT 79.290 64.640 79.610 65.840 ;
        RECT 76.090 63.440 78.330 63.840 ;
        RECT 79.930 63.280 80.890 67.170 ;
        RECT 74.170 63.040 75.150 63.280 ;
        RECT 79.930 63.040 80.910 63.280 ;
        RECT 0.470 55.740 26.850 56.300 ;
        RECT 0.470 55.190 5.300 55.740 ;
        RECT 0.470 54.630 26.750 55.190 ;
        RECT 0.470 38.710 5.300 54.630 ;
        RECT 6.290 52.670 7.730 53.870 ;
        RECT 7.370 49.070 7.730 52.670 ;
        RECT 8.450 52.670 9.890 53.870 ;
        RECT 8.450 49.070 8.810 52.670 ;
        RECT 9.530 49.070 9.890 52.670 ;
        RECT 10.610 52.670 12.050 53.870 ;
        RECT 10.610 49.070 10.970 52.670 ;
        RECT 11.690 49.070 12.050 52.670 ;
        RECT 12.770 52.670 14.210 53.870 ;
        RECT 12.770 49.070 13.130 52.670 ;
        RECT 13.850 49.070 14.210 52.670 ;
        RECT 14.930 52.670 16.370 53.870 ;
        RECT 14.930 49.070 15.290 52.670 ;
        RECT 16.010 49.070 16.370 52.670 ;
        RECT 17.090 52.670 18.530 53.870 ;
        RECT 17.090 49.070 17.450 52.670 ;
        RECT 18.170 49.070 18.530 52.670 ;
        RECT 19.250 52.670 20.690 53.870 ;
        RECT 19.250 49.070 19.610 52.670 ;
        RECT 20.330 49.070 20.690 52.670 ;
        RECT 21.410 52.670 22.850 53.870 ;
        RECT 21.410 49.070 21.770 52.670 ;
        RECT 22.490 49.070 22.850 52.670 ;
        RECT 23.570 52.670 25.010 53.870 ;
        RECT 23.570 49.070 23.930 52.670 ;
        RECT 7.370 39.470 8.810 41.870 ;
        RECT 9.530 39.470 10.970 41.870 ;
        RECT 11.690 39.470 13.130 41.870 ;
        RECT 13.850 39.470 15.290 41.870 ;
        RECT 16.010 39.470 17.450 41.870 ;
        RECT 18.170 39.470 19.610 41.870 ;
        RECT 20.330 39.470 21.770 41.870 ;
        RECT 22.490 39.470 23.930 41.870 ;
        RECT 26.190 38.710 26.750 54.630 ;
        RECT 29.020 48.400 29.980 58.170 ;
        RECT 30.940 55.900 33.180 56.300 ;
        RECT 30.300 53.900 30.620 55.100 ;
        RECT 31.580 54.300 33.820 54.700 ;
        RECT 34.140 53.900 34.460 55.100 ;
        RECT 30.940 52.700 33.180 53.100 ;
        RECT 30.940 51.790 33.180 52.190 ;
        RECT 30.300 49.790 30.620 50.990 ;
        RECT 31.580 50.190 33.820 50.590 ;
        RECT 34.140 49.790 34.460 50.990 ;
        RECT 30.940 48.590 33.180 48.990 ;
        RECT 34.780 48.400 35.740 58.100 ;
        RECT 38.930 48.440 39.890 58.100 ;
        RECT 40.850 55.940 43.090 56.340 ;
        RECT 40.210 53.940 40.530 55.140 ;
        RECT 41.490 54.340 43.730 54.740 ;
        RECT 44.050 53.940 44.370 55.140 ;
        RECT 40.850 52.740 43.090 53.140 ;
        RECT 40.850 51.830 43.090 52.230 ;
        RECT 40.210 49.830 40.530 51.030 ;
        RECT 41.490 50.230 43.730 50.630 ;
        RECT 44.050 49.830 44.370 51.030 ;
        RECT 40.850 48.630 43.090 49.030 ;
        RECT 44.690 48.440 45.650 58.170 ;
        RECT 54.550 54.060 55.510 60.230 ;
        RECT 56.470 57.660 58.710 58.060 ;
        RECT 55.830 55.660 56.150 56.860 ;
        RECT 57.110 56.060 59.350 56.460 ;
        RECT 59.670 55.660 59.990 56.860 ;
        RECT 56.470 54.460 58.710 54.860 ;
        RECT 60.310 54.060 61.270 60.290 ;
        RECT 63.060 57.770 64.020 61.490 ;
        RECT 64.980 61.100 67.220 61.500 ;
        RECT 68.810 61.490 69.780 61.900 ;
        RECT 64.340 59.100 64.660 60.300 ;
        RECT 65.620 59.500 67.860 59.900 ;
        RECT 68.180 59.100 68.500 60.300 ;
        RECT 64.980 57.900 67.220 58.300 ;
        RECT 68.820 57.770 69.780 61.490 ;
        RECT 74.190 58.880 75.150 63.040 ;
        RECT 76.110 62.480 78.350 62.880 ;
        RECT 75.470 60.480 75.790 61.680 ;
        RECT 76.750 60.880 78.990 61.280 ;
        RECT 79.310 60.480 79.630 61.680 ;
        RECT 76.110 59.280 78.350 59.680 ;
        RECT 79.950 58.880 80.910 63.040 ;
        RECT 83.540 58.880 84.500 65.020 ;
        RECT 85.460 62.480 87.700 62.880 ;
        RECT 84.820 60.480 85.140 61.680 ;
        RECT 86.100 60.880 88.340 61.280 ;
        RECT 88.660 60.480 88.980 61.680 ;
        RECT 85.460 59.280 87.700 59.680 ;
        RECT 89.300 58.880 90.260 64.990 ;
        RECT 63.050 57.500 64.020 57.770 ;
        RECT 68.810 57.500 69.780 57.770 ;
        RECT 29.010 48.190 29.980 48.400 ;
        RECT 34.770 48.190 35.740 48.400 ;
        RECT 38.920 48.230 39.890 48.440 ;
        RECT 44.680 48.230 45.650 48.440 ;
        RECT 54.800 52.610 59.300 52.650 ;
        RECT 63.050 52.610 64.010 57.500 ;
        RECT 64.970 56.970 67.210 57.370 ;
        RECT 64.330 54.970 64.650 56.170 ;
        RECT 65.610 55.370 67.850 55.770 ;
        RECT 68.170 54.970 68.490 56.170 ;
        RECT 64.970 53.770 67.210 54.170 ;
        RECT 68.810 52.660 69.770 57.500 ;
        RECT 74.120 52.660 75.080 57.760 ;
        RECT 76.040 56.960 78.280 57.360 ;
        RECT 75.400 54.960 75.720 56.160 ;
        RECT 76.680 55.360 78.920 55.760 ;
        RECT 79.240 54.960 79.560 56.160 ;
        RECT 76.040 53.760 78.280 54.160 ;
        RECT 76.040 52.660 77.000 53.210 ;
        RECT 79.880 52.660 80.840 57.760 ;
        RECT 64.930 52.610 80.840 52.660 ;
        RECT 54.800 51.860 80.840 52.610 ;
        RECT 54.800 50.360 81.190 51.860 ;
        RECT 92.580 50.360 93.780 76.150 ;
        RECT 149.810 76.140 159.340 76.150 ;
        RECT 138.410 71.670 139.470 73.750 ;
        RECT 138.380 70.510 139.470 71.670 ;
        RECT 138.380 69.350 139.440 70.510 ;
        RECT 138.050 69.330 139.440 69.350 ;
        RECT 107.000 68.920 129.200 69.240 ;
        RECT 136.130 69.230 142.880 69.330 ;
        RECT 105.470 68.680 129.200 68.920 ;
        RECT 105.470 52.760 107.560 68.680 ;
        RECT 108.740 66.720 110.180 67.920 ;
        RECT 109.820 63.120 110.180 66.720 ;
        RECT 110.900 66.720 112.340 67.920 ;
        RECT 110.900 63.120 111.260 66.720 ;
        RECT 111.980 63.120 112.340 66.720 ;
        RECT 113.060 66.720 114.500 67.920 ;
        RECT 113.060 63.120 113.420 66.720 ;
        RECT 114.140 63.120 114.500 66.720 ;
        RECT 115.220 66.720 116.660 67.920 ;
        RECT 115.220 63.120 115.580 66.720 ;
        RECT 116.300 63.120 116.660 66.720 ;
        RECT 117.380 66.720 118.820 67.920 ;
        RECT 117.380 63.120 117.740 66.720 ;
        RECT 118.460 63.120 118.820 66.720 ;
        RECT 119.540 66.720 120.980 67.920 ;
        RECT 119.540 63.120 119.900 66.720 ;
        RECT 120.620 63.120 120.980 66.720 ;
        RECT 121.700 66.720 123.140 67.920 ;
        RECT 121.700 63.120 122.060 66.720 ;
        RECT 122.780 63.120 123.140 66.720 ;
        RECT 123.860 66.720 125.300 67.920 ;
        RECT 123.860 63.120 124.220 66.720 ;
        RECT 124.940 63.120 125.300 66.720 ;
        RECT 126.020 66.720 127.460 67.920 ;
        RECT 126.020 63.120 126.380 66.720 ;
        RECT 109.820 53.520 111.260 55.920 ;
        RECT 111.980 53.520 113.420 55.920 ;
        RECT 114.140 53.520 115.580 55.920 ;
        RECT 116.300 53.520 117.740 55.920 ;
        RECT 118.460 53.520 119.900 55.920 ;
        RECT 120.620 53.520 122.060 55.920 ;
        RECT 122.780 53.520 124.220 55.920 ;
        RECT 124.940 53.520 126.380 55.920 ;
        RECT 128.640 52.760 129.200 68.680 ;
        RECT 136.120 68.370 142.880 69.230 ;
        RECT 136.120 68.270 142.850 68.370 ;
        RECT 136.130 65.230 137.090 68.270 ;
        RECT 138.050 65.370 139.010 68.270 ;
        RECT 141.890 65.230 142.850 68.270 ;
        RECT 136.120 64.080 137.090 65.230 ;
        RECT 138.040 64.430 140.280 64.830 ;
        RECT 136.120 61.320 137.080 64.080 ;
        RECT 141.880 63.850 142.850 65.230 ;
        RECT 137.400 62.430 137.720 63.630 ;
        RECT 138.680 62.830 140.920 63.230 ;
        RECT 141.240 62.430 141.560 63.630 ;
        RECT 136.120 60.830 137.110 61.320 ;
        RECT 138.040 61.230 140.280 61.630 ;
        RECT 141.880 61.600 142.840 63.850 ;
        RECT 141.880 60.830 142.870 61.600 ;
        RECT 136.150 60.210 137.110 60.830 ;
        RECT 141.910 60.210 142.870 60.830 ;
        RECT 136.140 58.480 137.110 60.210 ;
        RECT 138.060 59.410 140.300 59.810 ;
        RECT 136.140 55.810 137.100 58.480 ;
        RECT 137.420 57.410 137.740 58.610 ;
        RECT 138.700 57.810 140.940 58.210 ;
        RECT 141.260 57.410 141.580 58.610 ;
        RECT 141.900 58.500 142.870 60.210 ;
        RECT 138.060 56.210 140.300 56.610 ;
        RECT 141.900 55.810 142.860 58.500 ;
        RECT 105.470 52.200 129.200 52.760 ;
        RECT 105.470 51.650 107.560 52.200 ;
        RECT 105.470 51.090 129.100 51.650 ;
        RECT 105.470 51.080 107.560 51.090 ;
        RECT 54.800 49.800 94.080 50.360 ;
        RECT 54.800 49.780 81.190 49.800 ;
        RECT 29.010 39.890 29.970 48.190 ;
        RECT 30.930 47.600 33.170 48.000 ;
        RECT 30.290 45.600 30.610 46.800 ;
        RECT 31.570 46.000 33.810 46.400 ;
        RECT 34.130 45.600 34.450 46.800 ;
        RECT 30.930 44.400 33.170 44.800 ;
        RECT 30.930 43.490 33.170 43.890 ;
        RECT 30.290 41.490 30.610 42.690 ;
        RECT 31.570 41.890 33.810 42.290 ;
        RECT 34.130 41.490 34.450 42.690 ;
        RECT 30.930 40.290 33.170 40.690 ;
        RECT 34.770 39.890 35.730 48.190 ;
        RECT 38.920 39.930 39.880 48.230 ;
        RECT 40.840 47.640 43.080 48.040 ;
        RECT 40.200 45.640 40.520 46.840 ;
        RECT 41.480 46.040 43.720 46.440 ;
        RECT 44.040 45.640 44.360 46.840 ;
        RECT 40.840 44.440 43.080 44.840 ;
        RECT 40.840 43.530 43.080 43.930 ;
        RECT 40.200 41.530 40.520 42.730 ;
        RECT 41.480 41.930 43.720 42.330 ;
        RECT 44.040 41.530 44.360 42.730 ;
        RECT 40.840 40.330 43.080 40.730 ;
        RECT 44.680 39.930 45.640 48.230 ;
        RECT 0.470 38.150 26.750 38.710 ;
        RECT 0.470 37.720 5.300 38.150 ;
        RECT 0.470 37.160 26.690 37.720 ;
        RECT 0.470 21.240 5.300 37.160 ;
        RECT 6.230 35.200 7.670 36.400 ;
        RECT 7.310 31.600 7.670 35.200 ;
        RECT 8.390 35.200 9.830 36.400 ;
        RECT 8.390 31.600 8.750 35.200 ;
        RECT 9.470 31.600 9.830 35.200 ;
        RECT 10.550 35.200 11.990 36.400 ;
        RECT 10.550 31.600 10.910 35.200 ;
        RECT 11.630 31.600 11.990 35.200 ;
        RECT 12.710 35.200 14.150 36.400 ;
        RECT 12.710 31.600 13.070 35.200 ;
        RECT 13.790 31.600 14.150 35.200 ;
        RECT 14.870 35.200 16.310 36.400 ;
        RECT 14.870 31.600 15.230 35.200 ;
        RECT 15.950 31.600 16.310 35.200 ;
        RECT 17.030 35.200 18.470 36.400 ;
        RECT 17.030 31.600 17.390 35.200 ;
        RECT 18.110 31.600 18.470 35.200 ;
        RECT 19.190 35.200 20.630 36.400 ;
        RECT 19.190 31.600 19.550 35.200 ;
        RECT 20.270 31.600 20.630 35.200 ;
        RECT 21.350 35.200 22.790 36.400 ;
        RECT 21.350 31.600 21.710 35.200 ;
        RECT 22.430 31.600 22.790 35.200 ;
        RECT 23.510 35.200 24.950 36.400 ;
        RECT 23.510 31.600 23.870 35.200 ;
        RECT 7.310 22.000 8.750 24.400 ;
        RECT 9.470 22.000 10.910 24.400 ;
        RECT 11.630 22.000 13.070 24.400 ;
        RECT 13.790 22.000 15.230 24.400 ;
        RECT 15.950 22.000 17.390 24.400 ;
        RECT 18.110 22.000 19.550 24.400 ;
        RECT 20.270 22.000 21.710 24.400 ;
        RECT 22.430 22.000 23.870 24.400 ;
        RECT 26.130 21.240 26.690 37.160 ;
        RECT 29.020 29.540 29.980 36.530 ;
        RECT 30.940 35.730 33.180 36.130 ;
        RECT 30.300 33.730 30.620 34.930 ;
        RECT 31.580 34.130 33.820 34.530 ;
        RECT 34.140 33.730 34.460 34.930 ;
        RECT 30.940 32.530 33.180 32.930 ;
        RECT 30.940 29.540 31.900 31.420 ;
        RECT 34.780 29.540 35.740 36.530 ;
        RECT 38.940 29.540 39.900 36.520 ;
        RECT 40.860 35.720 43.100 36.120 ;
        RECT 40.220 33.720 40.540 34.920 ;
        RECT 41.500 34.120 43.740 34.520 ;
        RECT 44.060 33.720 44.380 34.920 ;
        RECT 40.860 32.520 43.100 32.920 ;
        RECT 40.860 29.540 41.820 31.540 ;
        RECT 44.700 29.540 45.660 36.520 ;
        RECT 29.020 29.530 45.660 29.540 ;
        RECT 0.470 20.830 26.690 21.240 ;
        RECT 28.860 28.560 45.660 29.530 ;
        RECT 28.860 20.830 45.210 28.560 ;
        RECT 54.800 25.920 59.300 49.780 ;
        RECT 65.960 45.180 66.920 45.230 ;
        RECT 62.140 44.220 66.920 45.180 ;
        RECT 60.200 38.730 61.160 43.990 ;
        RECT 62.120 42.050 64.360 42.450 ;
        RECT 61.480 40.050 61.800 41.250 ;
        RECT 62.760 40.450 65.000 40.850 ;
        RECT 65.320 40.050 65.640 41.250 ;
        RECT 62.120 38.850 64.360 39.250 ;
        RECT 65.960 38.730 66.920 44.220 ;
        RECT 60.200 38.450 61.170 38.730 ;
        RECT 65.960 38.450 66.930 38.730 ;
        RECT 60.210 34.330 61.170 38.450 ;
        RECT 62.130 37.930 64.370 38.330 ;
        RECT 61.490 35.930 61.810 37.130 ;
        RECT 62.770 36.330 65.010 36.730 ;
        RECT 65.330 35.930 65.650 37.130 ;
        RECT 62.130 34.730 64.370 35.130 ;
        RECT 65.970 34.330 66.930 38.450 ;
        RECT 70.750 33.960 71.310 49.780 ;
        RECT 71.820 47.920 73.930 49.120 ;
        RECT 73.570 44.320 73.930 47.920 ;
        RECT 74.650 47.920 76.090 49.120 ;
        RECT 74.650 44.320 75.010 47.920 ;
        RECT 75.730 44.320 76.090 47.920 ;
        RECT 76.810 47.920 78.890 49.120 ;
        RECT 76.810 44.320 77.170 47.920 ;
        RECT 73.570 34.720 75.010 37.120 ;
        RECT 75.730 34.720 77.170 37.120 ;
        RECT 79.430 33.960 79.990 49.780 ;
        RECT 70.750 33.860 79.990 33.960 ;
        RECT 80.520 33.880 81.080 49.780 ;
        RECT 81.540 49.040 83.410 49.110 ;
        RECT 81.540 47.910 83.700 49.040 ;
        RECT 82.260 47.840 83.700 47.910 ;
        RECT 83.340 44.240 83.700 47.840 ;
        RECT 84.420 47.840 85.860 49.040 ;
        RECT 84.420 44.240 84.780 47.840 ;
        RECT 85.500 44.240 85.860 47.840 ;
        RECT 86.580 47.840 88.020 49.040 ;
        RECT 86.580 44.240 86.940 47.840 ;
        RECT 87.660 44.240 88.020 47.840 ;
        RECT 88.740 47.840 90.180 49.040 ;
        RECT 88.740 44.240 89.100 47.840 ;
        RECT 89.820 44.240 90.180 47.840 ;
        RECT 90.900 47.840 92.850 49.040 ;
        RECT 90.900 44.240 91.260 47.840 ;
        RECT 83.340 34.640 84.780 37.040 ;
        RECT 85.500 34.640 86.940 37.040 ;
        RECT 87.660 34.640 89.100 37.040 ;
        RECT 89.820 34.640 91.260 37.040 ;
        RECT 93.520 33.880 94.080 49.800 ;
        RECT 80.520 33.860 94.080 33.880 ;
        RECT 70.750 33.400 94.080 33.860 ;
        RECT 70.830 33.320 94.080 33.400 ;
        RECT 105.470 35.170 107.460 51.080 ;
        RECT 108.640 49.130 110.080 50.330 ;
        RECT 109.720 45.530 110.080 49.130 ;
        RECT 110.800 49.130 112.240 50.330 ;
        RECT 110.800 45.530 111.160 49.130 ;
        RECT 111.880 45.530 112.240 49.130 ;
        RECT 112.960 49.130 114.400 50.330 ;
        RECT 112.960 45.530 113.320 49.130 ;
        RECT 114.040 45.530 114.400 49.130 ;
        RECT 115.120 49.130 116.560 50.330 ;
        RECT 115.120 45.530 115.480 49.130 ;
        RECT 116.200 45.530 116.560 49.130 ;
        RECT 117.280 49.130 118.720 50.330 ;
        RECT 117.280 45.530 117.640 49.130 ;
        RECT 118.360 45.530 118.720 49.130 ;
        RECT 119.440 49.130 120.880 50.330 ;
        RECT 119.440 45.530 119.800 49.130 ;
        RECT 120.520 45.530 120.880 49.130 ;
        RECT 121.600 49.130 123.040 50.330 ;
        RECT 121.600 45.530 121.960 49.130 ;
        RECT 122.680 45.530 123.040 49.130 ;
        RECT 123.760 49.130 125.200 50.330 ;
        RECT 123.760 45.530 124.120 49.130 ;
        RECT 124.840 45.530 125.200 49.130 ;
        RECT 125.920 49.130 127.360 50.330 ;
        RECT 125.920 45.530 126.280 49.130 ;
        RECT 109.720 35.930 111.160 38.330 ;
        RECT 111.880 35.930 113.320 38.330 ;
        RECT 114.040 35.930 115.480 38.330 ;
        RECT 116.200 35.930 117.640 38.330 ;
        RECT 118.360 35.930 119.800 38.330 ;
        RECT 120.520 35.930 121.960 38.330 ;
        RECT 122.680 35.930 124.120 38.330 ;
        RECT 124.840 35.930 126.280 38.330 ;
        RECT 128.540 35.170 129.100 51.090 ;
        RECT 131.370 44.860 132.330 54.630 ;
        RECT 133.290 52.360 135.530 52.760 ;
        RECT 132.650 50.360 132.970 51.560 ;
        RECT 133.930 50.760 136.170 51.160 ;
        RECT 136.490 50.360 136.810 51.560 ;
        RECT 133.290 49.160 135.530 49.560 ;
        RECT 133.290 48.250 135.530 48.650 ;
        RECT 132.650 46.250 132.970 47.450 ;
        RECT 133.930 46.650 136.170 47.050 ;
        RECT 136.490 46.250 136.810 47.450 ;
        RECT 133.290 45.050 135.530 45.450 ;
        RECT 137.130 44.860 138.090 54.560 ;
        RECT 141.280 44.900 142.240 54.560 ;
        RECT 143.200 52.400 145.440 52.800 ;
        RECT 142.560 50.400 142.880 51.600 ;
        RECT 143.840 50.800 146.080 51.200 ;
        RECT 146.400 50.400 146.720 51.600 ;
        RECT 143.200 49.200 145.440 49.600 ;
        RECT 143.200 48.290 145.440 48.690 ;
        RECT 142.560 46.290 142.880 47.490 ;
        RECT 143.840 46.690 146.080 47.090 ;
        RECT 146.400 46.290 146.720 47.490 ;
        RECT 143.200 45.090 145.440 45.490 ;
        RECT 147.040 44.900 148.000 54.630 ;
        RECT 131.360 44.650 132.330 44.860 ;
        RECT 137.120 44.650 138.090 44.860 ;
        RECT 141.270 44.690 142.240 44.900 ;
        RECT 147.030 44.690 148.000 44.900 ;
        RECT 131.360 36.350 132.320 44.650 ;
        RECT 133.280 44.060 135.520 44.460 ;
        RECT 132.640 42.060 132.960 43.260 ;
        RECT 133.920 42.460 136.160 42.860 ;
        RECT 136.480 42.060 136.800 43.260 ;
        RECT 133.280 40.860 135.520 41.260 ;
        RECT 133.280 39.950 135.520 40.350 ;
        RECT 132.640 37.950 132.960 39.150 ;
        RECT 133.920 38.350 136.160 38.750 ;
        RECT 136.480 37.950 136.800 39.150 ;
        RECT 133.280 36.750 135.520 37.150 ;
        RECT 137.120 36.350 138.080 44.650 ;
        RECT 141.270 36.390 142.230 44.690 ;
        RECT 143.190 44.100 145.430 44.500 ;
        RECT 142.550 42.100 142.870 43.300 ;
        RECT 143.830 42.500 146.070 42.900 ;
        RECT 146.390 42.100 146.710 43.300 ;
        RECT 143.190 40.900 145.430 41.300 ;
        RECT 143.190 39.990 145.430 40.390 ;
        RECT 142.550 37.990 142.870 39.190 ;
        RECT 143.830 38.390 146.070 38.790 ;
        RECT 146.390 37.990 146.710 39.190 ;
        RECT 143.190 36.790 145.430 37.190 ;
        RECT 147.030 36.390 147.990 44.690 ;
        RECT 105.470 34.610 129.100 35.170 ;
        RECT 105.470 34.180 107.460 34.610 ;
        RECT 105.470 33.620 129.040 34.180 ;
        RECT 0.470 20.655 45.210 20.830 ;
        RECT 48.420 24.745 59.300 25.920 ;
        RECT 48.420 20.655 49.595 24.745 ;
        RECT 49.905 20.965 53.375 24.435 ;
        RECT 53.685 20.655 59.300 24.745 ;
        RECT 62.200 32.600 66.240 32.930 ;
        RECT 70.830 32.600 92.960 33.320 ;
        RECT 62.200 32.140 92.960 32.600 ;
        RECT 62.200 32.105 93.060 32.140 ;
        RECT 62.200 31.785 66.340 32.105 ;
        RECT 70.720 31.990 93.060 32.105 ;
        RECT 70.720 31.785 72.870 31.990 ;
        RECT 77.330 31.785 78.360 31.990 ;
        RECT 62.200 31.425 78.360 31.785 ;
        RECT 62.200 27.335 66.375 31.425 ;
        RECT 66.685 27.645 70.155 31.115 ;
        RECT 70.465 27.335 73.095 31.425 ;
        RECT 73.405 27.645 76.875 31.115 ;
        RECT 77.185 27.335 78.360 31.425 ;
        RECT 62.200 26.975 78.360 27.335 ;
        RECT 62.200 26.655 66.340 26.975 ;
        RECT 70.720 26.655 72.870 26.975 ;
        RECT 77.330 26.655 78.360 26.975 ;
        RECT 62.200 26.390 78.360 26.655 ;
        RECT 78.700 31.775 79.610 31.990 ;
        RECT 84.090 31.775 86.350 31.990 ;
        RECT 78.700 31.765 86.350 31.775 ;
        RECT 78.700 31.415 91.065 31.765 ;
        RECT 78.700 27.325 79.875 31.415 ;
        RECT 83.965 31.405 91.065 31.415 ;
        RECT 80.185 27.635 83.655 31.105 ;
        RECT 83.965 27.325 86.615 31.405 ;
        RECT 86.925 27.625 90.395 31.095 ;
        RECT 78.700 27.315 86.615 27.325 ;
        RECT 90.705 27.315 91.065 31.405 ;
        RECT 78.700 26.965 91.065 27.315 ;
        RECT 78.700 26.645 79.610 26.965 ;
        RECT 84.090 26.955 91.065 26.965 ;
        RECT 84.090 26.645 86.350 26.955 ;
        RECT 78.700 26.635 86.350 26.645 ;
        RECT 91.385 26.635 93.060 31.990 ;
        RECT 78.700 26.390 93.060 26.635 ;
        RECT 62.200 25.300 93.060 26.390 ;
        RECT 62.200 25.205 78.380 25.300 ;
        RECT 62.200 24.885 66.340 25.205 ;
        RECT 70.720 24.885 72.870 25.205 ;
        RECT 77.330 24.885 78.380 25.205 ;
        RECT 62.200 24.525 78.380 24.885 ;
        RECT 62.200 20.655 66.375 24.525 ;
        RECT 66.685 20.745 70.155 24.215 ;
        RECT 0.470 20.435 66.375 20.655 ;
        RECT 70.465 20.435 73.115 24.525 ;
        RECT 73.425 20.745 76.895 24.215 ;
        RECT 77.205 20.435 78.380 24.525 ;
        RECT 0.470 20.110 78.380 20.435 ;
        RECT 78.690 25.205 93.060 25.300 ;
        RECT 78.690 24.885 79.610 25.205 ;
        RECT 84.090 24.885 86.350 25.205 ;
        RECT 78.690 24.525 91.055 24.885 ;
        RECT 78.690 20.435 79.865 24.525 ;
        RECT 80.175 20.745 83.645 24.215 ;
        RECT 83.955 20.435 86.605 24.525 ;
        RECT 86.915 20.745 90.385 24.215 ;
        RECT 90.695 20.435 91.055 24.525 ;
        RECT 78.690 20.110 91.055 20.435 ;
        RECT 91.375 20.110 93.060 25.205 ;
        RECT 0.470 19.530 93.060 20.110 ;
        RECT 0.470 17.790 93.540 19.530 ;
        RECT 95.600 17.790 96.560 26.350 ;
        RECT 97.520 24.750 99.120 25.150 ;
        RECT 96.880 23.550 97.200 24.750 ;
        RECT 98.160 23.950 99.760 24.350 ;
        RECT 100.080 23.550 100.400 24.750 ;
        RECT 97.520 23.150 99.120 23.550 ;
        RECT 97.640 17.790 98.480 21.410 ;
        RECT 100.720 17.790 101.680 26.350 ;
        RECT 103.040 17.790 104.360 19.920 ;
        RECT 105.470 17.790 107.460 33.620 ;
        RECT 108.580 31.660 110.020 32.860 ;
        RECT 109.660 28.060 110.020 31.660 ;
        RECT 110.740 31.660 112.180 32.860 ;
        RECT 110.740 28.060 111.100 31.660 ;
        RECT 111.820 28.060 112.180 31.660 ;
        RECT 112.900 31.660 114.340 32.860 ;
        RECT 112.900 28.060 113.260 31.660 ;
        RECT 113.980 28.060 114.340 31.660 ;
        RECT 115.060 31.660 116.500 32.860 ;
        RECT 115.060 28.060 115.420 31.660 ;
        RECT 116.140 28.060 116.500 31.660 ;
        RECT 117.220 31.660 118.660 32.860 ;
        RECT 117.220 28.060 117.580 31.660 ;
        RECT 118.300 28.060 118.660 31.660 ;
        RECT 119.380 31.660 120.820 32.860 ;
        RECT 119.380 28.060 119.740 31.660 ;
        RECT 120.460 28.060 120.820 31.660 ;
        RECT 121.540 31.660 122.980 32.860 ;
        RECT 121.540 28.060 121.900 31.660 ;
        RECT 122.620 28.060 122.980 31.660 ;
        RECT 123.700 31.660 125.140 32.860 ;
        RECT 123.700 28.060 124.060 31.660 ;
        RECT 124.780 28.060 125.140 31.660 ;
        RECT 125.860 31.660 127.300 32.860 ;
        RECT 125.860 28.060 126.220 31.660 ;
        RECT 109.660 18.460 111.100 20.860 ;
        RECT 111.820 18.460 113.260 20.860 ;
        RECT 113.980 18.460 115.420 20.860 ;
        RECT 116.140 18.460 117.580 20.860 ;
        RECT 118.300 18.460 119.740 20.860 ;
        RECT 120.460 18.460 121.900 20.860 ;
        RECT 122.620 18.460 124.060 20.860 ;
        RECT 124.780 18.460 126.220 20.860 ;
        RECT 128.480 17.790 129.040 33.620 ;
        RECT 131.370 26.000 132.330 32.990 ;
        RECT 133.290 32.190 135.530 32.590 ;
        RECT 132.650 30.190 132.970 31.390 ;
        RECT 133.930 30.590 136.170 30.990 ;
        RECT 136.490 30.190 136.810 31.390 ;
        RECT 133.290 28.990 135.530 29.390 ;
        RECT 133.290 26.000 134.250 27.880 ;
        RECT 137.130 26.000 138.090 32.990 ;
        RECT 141.290 26.000 142.250 32.980 ;
        RECT 143.210 32.180 145.450 32.580 ;
        RECT 142.570 30.180 142.890 31.380 ;
        RECT 143.850 30.580 146.090 30.980 ;
        RECT 146.410 30.180 146.730 31.380 ;
        RECT 143.210 28.980 145.450 29.380 ;
        RECT 143.210 26.000 144.170 28.000 ;
        RECT 147.050 26.000 148.010 32.980 ;
        RECT 131.370 25.990 148.010 26.000 ;
        RECT 131.210 25.970 148.010 25.990 ;
        RECT 150.730 25.970 159.300 76.140 ;
        RECT 131.210 19.250 159.300 25.970 ;
        RECT 131.210 17.790 159.280 19.250 ;
        RECT 0.470 6.990 159.280 17.790 ;
        RECT 0.470 6.830 153.180 6.990 ;
        RECT 0.500 6.550 153.180 6.830 ;
        RECT 0.500 6.480 4.530 6.550 ;
      LAYER met1 ;
        RECT 12.520 211.990 108.520 212.390 ;
        RECT 12.520 211.870 108.620 211.990 ;
        RECT 12.380 210.390 108.620 211.870 ;
        RECT 11.740 189.870 12.060 209.330 ;
        RECT 12.380 191.230 13.340 210.390 ;
        RECT 14.300 189.870 15.260 209.330 ;
        RECT 20.740 189.870 21.060 208.830 ;
        RECT 21.380 191.230 22.340 210.390 ;
        RECT 23.300 205.880 24.260 208.830 ;
        RECT 23.290 193.860 24.270 205.880 ;
        RECT 23.300 189.870 24.260 193.860 ;
        RECT 29.740 189.870 30.060 208.830 ;
        RECT 30.380 191.230 31.340 210.390 ;
        RECT 32.300 189.870 33.260 208.830 ;
        RECT 38.740 189.870 39.060 208.830 ;
        RECT 39.380 191.230 40.340 210.390 ;
        RECT 41.300 189.870 42.260 208.830 ;
        RECT 47.740 201.710 48.060 201.830 ;
        RECT 47.420 189.870 48.060 201.710 ;
        RECT 48.380 198.230 49.340 210.390 ;
        RECT 11.540 189.230 48.060 189.870 ;
        RECT 11.540 188.910 48.000 189.230 ;
        RECT 32.360 187.290 33.560 188.910 ;
        RECT 50.300 187.930 51.260 201.830 ;
        RECT 56.740 189.050 57.060 208.830 ;
        RECT 57.380 191.230 58.340 210.390 ;
        RECT 59.300 204.370 60.260 208.830 ;
        RECT 59.270 203.410 60.290 204.370 ;
        RECT 59.300 195.880 60.260 201.830 ;
        RECT 49.570 187.870 51.260 187.930 ;
        RECT 53.860 188.730 57.060 189.050 ;
        RECT 59.300 188.880 60.260 194.830 ;
        RECT 13.420 185.890 16.120 187.290 ;
        RECT 32.220 185.890 33.720 187.290 ;
        RECT 39.380 186.910 51.300 187.870 ;
        RECT 13.420 169.290 14.620 185.890 ;
        RECT 38.740 175.230 39.060 186.580 ;
        RECT 39.380 175.230 40.340 186.910 ;
        RECT 41.300 173.870 42.260 186.330 ;
        RECT 47.740 175.230 48.060 186.580 ;
        RECT 48.380 175.230 49.340 186.910 ;
        RECT 49.570 186.850 50.530 186.910 ;
        RECT 38.540 172.910 48.500 173.870 ;
        RECT 50.300 173.550 51.260 185.830 ;
        RECT 53.860 173.550 54.180 188.730 ;
        RECT 50.300 173.030 54.180 173.550 ;
        RECT 13.420 167.890 16.120 169.290 ;
        RECT 38.740 162.230 39.060 172.910 ;
        RECT 39.380 161.860 40.340 170.830 ;
        RECT 41.300 162.230 42.260 172.910 ;
        RECT 47.740 162.230 48.060 172.910 ;
        RECT 44.510 161.870 45.470 161.930 ;
        RECT 48.380 161.870 49.340 170.830 ;
        RECT 50.300 162.230 51.260 173.030 ;
        RECT 53.860 166.550 54.180 173.030 ;
        RECT 53.860 166.230 56.210 166.550 ;
        RECT 43.600 161.860 49.340 161.870 ;
        RECT 39.380 160.920 49.340 161.860 ;
        RECT 39.380 160.910 40.340 160.920 ;
        RECT 43.600 160.910 49.340 160.920 ;
        RECT 44.510 160.850 45.470 160.910 ;
        RECT 35.890 159.050 37.150 160.250 ;
        RECT 61.520 159.670 63.520 210.390 ;
        RECT 66.780 187.930 67.740 201.830 ;
        RECT 68.700 198.230 69.660 210.390 ;
        RECT 69.980 201.710 70.300 201.830 ;
        RECT 69.980 189.870 70.620 201.710 ;
        RECT 75.780 189.870 76.740 208.830 ;
        RECT 77.700 191.230 78.660 210.390 ;
        RECT 78.980 189.870 79.300 208.830 ;
        RECT 84.780 189.870 85.740 208.830 ;
        RECT 86.700 191.230 87.660 210.390 ;
        RECT 87.980 189.870 88.300 208.830 ;
        RECT 93.780 205.880 94.740 208.830 ;
        RECT 93.770 193.860 94.750 205.880 ;
        RECT 93.780 189.870 94.740 193.860 ;
        RECT 95.700 191.230 96.660 210.390 ;
        RECT 96.980 189.870 97.300 208.830 ;
        RECT 102.780 189.870 103.740 209.330 ;
        RECT 104.700 191.230 105.660 210.390 ;
        RECT 107.420 210.190 108.620 210.390 ;
        RECT 110.720 210.190 112.120 210.290 ;
        RECT 105.980 189.870 106.300 209.330 ;
        RECT 107.420 208.990 112.120 210.190 ;
        RECT 110.720 208.890 112.120 208.990 ;
        RECT 115.320 208.890 117.620 210.290 ;
        RECT 116.420 192.290 117.620 208.890 ;
        RECT 109.920 190.890 112.120 192.290 ;
        RECT 115.320 190.890 117.620 192.290 ;
        RECT 69.980 189.230 106.500 189.870 ;
        RECT 70.040 188.910 106.500 189.230 ;
        RECT 66.780 187.870 68.470 187.930 ;
        RECT 66.740 186.910 78.660 187.870 ;
        RECT 84.480 187.290 85.680 188.910 ;
        RECT 67.510 186.850 68.470 186.910 ;
        RECT 66.780 173.440 67.740 185.830 ;
        RECT 68.700 175.230 69.660 186.910 ;
        RECT 69.980 175.230 70.300 186.580 ;
        RECT 75.780 173.870 76.740 186.330 ;
        RECT 77.700 175.230 78.660 186.910 ;
        RECT 78.980 175.230 79.300 186.580 ;
        RECT 84.320 185.890 85.820 187.290 ;
        RECT 101.920 185.890 104.620 187.290 ;
        RECT 64.270 173.140 67.740 173.440 ;
        RECT 64.270 160.340 64.570 173.140 ;
        RECT 66.780 162.230 67.740 173.140 ;
        RECT 69.540 172.910 79.500 173.870 ;
        RECT 68.700 161.870 69.660 170.830 ;
        RECT 69.980 162.230 70.300 172.910 ;
        RECT 75.780 162.230 76.740 172.910 ;
        RECT 72.570 161.870 73.530 161.930 ;
        RECT 68.700 161.860 74.440 161.870 ;
        RECT 77.700 161.860 78.660 170.830 ;
        RECT 78.980 162.230 79.300 172.910 ;
        RECT 103.420 169.290 104.620 185.890 ;
        RECT 109.920 174.250 111.120 190.890 ;
        RECT 116.600 174.250 117.620 176.230 ;
        RECT 109.920 172.990 112.010 174.250 ;
        RECT 110.810 172.930 112.010 172.990 ;
        RECT 115.430 172.930 117.620 174.250 ;
        RECT 101.920 167.890 104.620 169.290 ;
        RECT 68.700 160.920 78.660 161.860 ;
        RECT 68.700 160.910 74.440 160.920 ;
        RECT 77.700 160.910 78.660 160.920 ;
        RECT 72.570 160.850 73.530 160.910 ;
        RECT 64.270 160.040 72.600 160.340 ;
        RECT 13.920 149.890 16.120 151.290 ;
        RECT 32.390 151.190 33.590 151.250 ;
        RECT 35.920 151.190 37.120 159.050 ;
        RECT 61.520 158.710 65.830 159.670 ;
        RECT 51.170 158.440 51.470 158.470 ;
        RECT 49.940 158.140 51.470 158.440 ;
        RECT 51.170 158.110 51.470 158.140 ;
        RECT 32.390 149.990 37.120 151.190 ;
        RECT 39.620 153.090 59.120 156.490 ;
        RECT 61.520 156.390 63.520 158.710 ;
        RECT 65.940 156.010 66.240 158.600 ;
        RECT 66.740 157.440 67.620 157.780 ;
        RECT 69.440 157.440 70.320 157.780 ;
        RECT 72.300 156.980 72.600 160.040 ;
        RECT 71.080 156.330 71.960 156.360 ;
        RECT 71.080 155.450 75.190 156.330 ;
        RECT 116.420 156.250 117.620 172.930 ;
        RECT 71.080 155.420 71.960 155.450 ;
        RECT 115.430 154.990 117.620 156.250 ;
        RECT 115.430 154.930 116.630 154.990 ;
        RECT 67.840 154.040 68.140 154.100 ;
        RECT 65.340 153.740 68.140 154.040 ;
        RECT 67.840 153.680 68.140 153.740 ;
        RECT 68.620 153.440 69.500 153.480 ;
        RECT 68.620 153.140 70.120 153.440 ;
        RECT 32.390 149.930 33.590 149.990 ;
        RECT 13.920 133.290 15.120 149.890 ;
        RECT 39.620 140.390 43.020 153.090 ;
        RECT 48.920 148.265 50.120 151.020 ;
        RECT 47.845 145.215 50.895 148.265 ;
        RECT 55.820 140.390 59.120 153.090 ;
        RECT 65.920 152.340 66.800 152.680 ;
        RECT 68.620 152.340 69.500 152.680 ;
        RECT 65.920 151.840 66.800 151.880 ;
        RECT 65.920 151.540 67.420 151.840 ;
        RECT 64.120 151.140 65.000 151.480 ;
        RECT 64.120 149.840 65.000 149.880 ;
        RECT 39.620 137.090 59.120 140.390 ;
        RECT 63.520 149.540 65.000 149.840 ;
        RECT 63.520 137.840 63.820 149.540 ;
        RECT 65.920 149.140 66.800 149.480 ;
        RECT 65.920 148.640 66.800 148.680 ;
        RECT 67.120 148.640 67.420 151.540 ;
        RECT 69.820 150.640 70.120 153.140 ;
        RECT 102.890 152.490 104.090 152.550 ;
        RECT 100.890 151.290 104.090 152.490 ;
        RECT 102.890 151.230 104.090 151.290 ;
        RECT 70.420 150.640 71.300 150.680 ;
        RECT 69.820 150.340 71.300 150.640 ;
        RECT 68.620 149.940 69.500 150.280 ;
        RECT 65.920 148.340 67.420 148.640 ;
        RECT 70.420 148.240 71.300 148.280 ;
        RECT 70.420 147.940 71.920 148.240 ;
        RECT 70.420 147.440 71.300 147.480 ;
        RECT 69.820 147.140 71.300 147.440 ;
        RECT 65.920 146.740 66.800 147.080 ;
        RECT 68.620 146.740 69.500 147.080 ;
        RECT 68.620 146.240 69.500 146.280 ;
        RECT 69.820 146.240 70.120 147.140 ;
        RECT 68.620 145.940 70.120 146.240 ;
        RECT 64.120 145.840 65.000 145.880 ;
        RECT 64.120 145.540 65.620 145.840 ;
        RECT 65.320 144.640 65.620 145.540 ;
        RECT 65.920 145.140 66.800 145.480 ;
        RECT 68.620 145.140 69.500 145.480 ;
        RECT 65.920 144.640 66.800 144.680 ;
        RECT 65.320 144.340 66.800 144.640 ;
        RECT 69.820 143.440 70.120 145.940 ;
        RECT 70.420 144.240 71.300 144.280 ;
        RECT 71.620 144.240 71.920 147.940 ;
        RECT 70.420 143.940 71.920 144.240 ;
        RECT 70.420 143.440 71.300 143.480 ;
        RECT 69.820 143.140 71.300 143.440 ;
        RECT 65.920 142.740 66.800 143.080 ;
        RECT 68.620 142.740 69.500 143.080 ;
        RECT 64.120 141.840 65.000 141.880 ;
        RECT 64.120 141.540 65.020 141.840 ;
        RECT 64.720 141.240 65.620 141.540 ;
        RECT 65.320 138.240 65.620 141.240 ;
        RECT 65.920 140.340 66.800 140.680 ;
        RECT 68.620 140.340 69.500 140.680 ;
        RECT 70.810 140.210 71.230 140.510 ;
        RECT 70.870 139.710 71.170 140.210 ;
        RECT 65.920 138.740 66.800 139.080 ;
        RECT 68.620 138.740 69.500 139.080 ;
        RECT 65.920 138.240 66.800 138.280 ;
        RECT 65.320 137.940 66.800 138.240 ;
        RECT 68.620 137.940 69.500 138.280 ;
        RECT 64.120 137.840 65.000 137.880 ;
        RECT 63.520 137.540 65.000 137.840 ;
        RECT 56.360 133.290 57.560 137.090 ;
        RECT 63.520 134.140 63.820 137.540 ;
        RECT 68.620 137.440 69.500 137.480 ;
        RECT 71.620 137.440 71.920 143.940 ;
        RECT 68.620 137.140 71.920 137.440 ;
        RECT 65.920 136.340 66.800 136.680 ;
        RECT 68.620 136.340 69.500 136.680 ;
        RECT 65.920 135.540 66.800 135.880 ;
        RECT 68.620 135.540 69.500 135.880 ;
        RECT 65.920 134.740 66.800 135.080 ;
        RECT 68.620 134.740 69.500 135.080 ;
        RECT 63.520 133.840 70.000 134.140 ;
        RECT 13.920 131.890 16.220 133.290 ;
        RECT 32.320 133.190 33.620 133.290 ;
        RECT 38.720 133.190 40.120 133.290 ;
        RECT 32.320 131.990 40.120 133.190 ;
        RECT 32.320 131.890 33.620 131.990 ;
        RECT 38.720 131.890 40.120 131.990 ;
        RECT 56.320 131.890 57.620 133.290 ;
        RECT 61.170 132.740 61.620 133.190 ;
        RECT 61.240 124.730 61.560 132.740 ;
        RECT 61.880 123.380 62.840 133.130 ;
        RECT 63.160 132.170 67.430 133.130 ;
        RECT 63.160 124.730 64.120 132.170 ;
        RECT 66.700 129.140 67.640 130.020 ;
        RECT 66.730 127.610 67.610 129.140 ;
        RECT 0.620 102.380 154.510 113.540 ;
        RECT 0.680 74.540 53.810 102.380 ;
        RECT 74.180 101.630 75.140 102.380 ;
        RECT 74.120 100.670 75.200 101.630 ;
        RECT 75.460 98.110 75.780 99.930 ;
        RECT 75.460 96.330 75.790 98.110 ;
        RECT 75.470 95.770 75.790 96.330 ;
        RECT 76.100 95.770 77.060 102.380 ;
        RECT 79.940 101.630 80.900 102.380 ;
        RECT 79.880 100.670 80.960 101.630 ;
        RECT 83.540 100.230 89.780 102.380 ;
        RECT 112.920 100.390 114.120 100.450 ;
        RECT 108.970 100.370 114.120 100.390 ;
        RECT 102.300 100.310 103.500 100.370 ;
        RECT 91.650 100.230 92.850 100.290 ;
        RECT 78.020 98.980 78.980 99.930 ;
        RECT 83.520 99.030 92.850 100.230 ;
        RECT 78.020 96.330 78.990 98.980 ;
        RECT 78.030 95.770 78.990 96.330 ;
        RECT 64.300 89.880 64.620 94.010 ;
        RECT 64.940 93.930 65.900 94.010 ;
        RECT 64.940 90.410 65.930 93.930 ;
        RECT 66.860 93.110 67.820 94.010 ;
        RECT 66.860 90.410 67.850 93.110 ;
        RECT 75.440 92.170 75.790 95.770 ;
        RECT 76.080 92.170 77.060 95.770 ;
        RECT 78.000 92.170 78.990 95.770 ;
        RECT 64.970 89.880 65.930 90.410 ;
        RECT 66.890 89.880 67.850 90.410 ;
        RECT 64.290 86.280 64.620 89.880 ;
        RECT 64.930 86.280 65.930 89.880 ;
        RECT 66.850 86.280 67.850 89.880 ;
        RECT 75.470 91.780 75.790 92.170 ;
        RECT 76.100 91.780 77.060 92.170 ;
        RECT 78.030 91.780 78.990 92.170 ;
        RECT 75.470 88.180 75.800 91.780 ;
        RECT 76.100 88.180 77.080 91.780 ;
        RECT 78.030 88.180 79.000 91.780 ;
        RECT 75.470 87.620 75.790 88.180 ;
        RECT 76.100 87.620 77.060 88.180 ;
        RECT 78.030 87.620 78.990 88.180 ;
        RECT 64.300 85.880 64.620 86.280 ;
        RECT 64.970 85.880 65.930 86.280 ;
        RECT 66.890 85.880 67.850 86.280 ;
        RECT 64.300 82.280 64.640 85.880 ;
        RECT 64.960 82.280 65.930 85.880 ;
        RECT 66.880 82.280 67.850 85.880 ;
        RECT 75.440 84.020 75.790 87.620 ;
        RECT 76.080 84.020 77.060 87.620 ;
        RECT 78.000 84.020 78.990 87.620 ;
        RECT 75.470 83.620 75.790 84.020 ;
        RECT 64.300 81.750 64.620 82.280 ;
        RECT 64.970 81.750 65.930 82.280 ;
        RECT 66.890 81.750 67.850 82.280 ;
        RECT 64.300 78.150 64.630 81.750 ;
        RECT 64.950 78.150 65.930 81.750 ;
        RECT 66.870 78.150 67.850 81.750 ;
        RECT 75.460 80.020 75.790 83.620 ;
        RECT 75.470 79.460 75.790 80.020 ;
        RECT 76.100 79.460 77.060 84.020 ;
        RECT 78.030 83.620 78.990 84.020 ;
        RECT 78.020 80.020 78.990 83.620 ;
        RECT 78.030 79.460 78.990 80.020 ;
        RECT 64.300 77.760 64.620 78.150 ;
        RECT 64.970 77.760 65.930 78.150 ;
        RECT 66.890 77.760 67.850 78.150 ;
        RECT 39.570 72.930 53.770 74.540 ;
        RECT 39.290 71.810 53.770 72.930 ;
        RECT 39.290 71.750 40.350 71.810 ;
        RECT 23.940 71.460 25.140 71.520 ;
        RECT 37.620 71.460 38.580 71.470 ;
        RECT 6.330 70.230 7.650 71.430 ;
        RECT 23.940 70.260 38.580 71.460 ;
        RECT 6.390 58.790 7.590 70.230 ;
        RECT 23.940 70.200 25.140 70.260 ;
        RECT 35.060 68.370 35.380 70.260 ;
        RECT 35.700 68.370 36.660 69.900 ;
        RECT 37.620 68.370 38.580 70.260 ;
        RECT 35.050 67.630 35.380 68.370 ;
        RECT 35.050 65.240 35.370 67.630 ;
        RECT 35.690 66.700 36.660 68.370 ;
        RECT 37.610 67.060 38.580 68.370 ;
        RECT 35.690 65.690 36.650 66.700 ;
        RECT 35.050 64.770 35.400 65.240 ;
        RECT 35.690 64.770 36.680 65.690 ;
        RECT 37.610 64.770 38.570 67.060 ;
        RECT 35.080 63.350 35.400 64.770 ;
        RECT 35.720 63.350 36.680 64.770 ;
        RECT 46.440 63.880 53.770 71.810 ;
        RECT 64.300 74.160 64.640 77.760 ;
        RECT 64.960 74.160 65.930 77.760 ;
        RECT 66.880 74.160 67.850 77.760 ;
        RECT 75.440 75.860 75.790 79.460 ;
        RECT 76.080 75.860 77.060 79.460 ;
        RECT 78.000 75.860 78.990 79.460 ;
        RECT 75.470 75.330 75.790 75.860 ;
        RECT 64.300 73.630 64.620 74.160 ;
        RECT 64.970 73.630 65.930 74.160 ;
        RECT 66.890 73.630 67.850 74.160 ;
        RECT 64.300 70.030 64.630 73.630 ;
        RECT 64.950 70.030 65.930 73.630 ;
        RECT 66.870 70.030 67.850 73.630 ;
        RECT 75.460 71.730 75.790 75.330 ;
        RECT 64.300 69.620 64.620 70.030 ;
        RECT 64.970 69.620 65.930 70.030 ;
        RECT 66.890 69.620 67.850 70.030 ;
        RECT 64.300 66.020 64.660 69.620 ;
        RECT 64.970 66.020 65.940 69.620 ;
        RECT 66.890 66.020 67.860 69.620 ;
        RECT 75.470 67.040 75.790 71.730 ;
        RECT 76.100 71.170 77.060 75.860 ;
        RECT 78.030 75.330 78.990 75.860 ;
        RECT 78.020 71.730 78.990 75.330 ;
        RECT 76.100 67.570 77.070 71.170 ;
        RECT 76.100 67.040 77.060 67.570 ;
        RECT 78.030 67.040 78.990 71.730 ;
        RECT 64.300 65.490 64.620 66.020 ;
        RECT 35.070 62.120 35.400 63.350 ;
        RECT 35.070 59.750 35.390 62.120 ;
        RECT 35.710 61.240 36.680 63.350 ;
        RECT 35.710 59.750 36.670 61.240 ;
        RECT 37.630 60.210 38.590 63.350 ;
        RECT 46.370 60.350 61.100 63.880 ;
        RECT 64.300 61.890 64.650 65.490 ;
        RECT 64.300 61.500 64.620 61.890 ;
        RECT 64.970 61.500 65.930 66.020 ;
        RECT 66.890 61.500 67.850 66.020 ;
        RECT 75.450 63.440 75.790 67.040 ;
        RECT 76.090 63.440 77.060 67.040 ;
        RECT 78.010 63.440 78.990 67.040 ;
        RECT 83.540 66.330 89.780 99.030 ;
        RECT 91.650 98.970 92.850 99.030 ;
        RECT 97.420 100.230 98.620 100.290 ;
        RECT 99.320 100.230 103.500 100.310 ;
        RECT 97.420 99.110 103.500 100.230 ;
        RECT 97.420 99.030 101.280 99.110 ;
        RECT 102.300 99.050 103.500 99.110 ;
        RECT 108.200 99.190 114.120 100.370 ;
        RECT 108.200 99.110 112.260 99.190 ;
        RECT 112.920 99.130 114.120 99.190 ;
        RECT 118.820 100.390 120.020 100.450 ;
        RECT 118.820 99.190 122.820 100.390 ;
        RECT 118.820 99.130 120.020 99.190 ;
        RECT 108.200 99.050 109.400 99.110 ;
        RECT 97.420 98.970 98.620 99.030 ;
        RECT 111.005 81.305 111.335 99.110 ;
        RECT 121.620 84.350 122.820 99.190 ;
        RECT 121.590 83.150 122.850 84.350 ;
        RECT 110.975 80.975 111.365 81.305 ;
        RECT 135.070 72.690 139.550 102.380 ;
        RECT 138.410 72.660 139.470 72.690 ;
        RECT 126.290 67.920 127.490 67.980 ;
        RECT 139.970 67.920 140.930 67.930 ;
        RECT 108.680 66.690 110.000 67.890 ;
        RECT 126.290 66.720 140.930 67.920 ;
        RECT 83.510 65.370 90.260 66.330 ;
        RECT 83.510 65.050 84.500 65.370 ;
        RECT 83.480 64.090 84.560 65.050 ;
        RECT 37.630 59.750 38.600 60.210 ;
        RECT 6.390 57.590 24.950 58.790 ;
        RECT 6.260 46.590 7.460 53.930 ;
        RECT 23.750 52.640 24.950 57.590 ;
        RECT 28.960 58.150 32.470 58.200 ;
        RECT 37.640 58.150 38.600 59.750 ;
        RECT 46.370 59.290 61.240 60.350 ;
        RECT 44.660 58.170 45.620 58.230 ;
        RECT 40.140 58.150 45.620 58.170 ;
        RECT 28.960 57.240 45.620 58.150 ;
        RECT 30.940 57.210 45.620 57.240 ;
        RECT 30.940 57.190 41.840 57.210 ;
        RECT 27.645 48.000 27.975 48.030 ;
        RECT 30.300 48.000 30.620 56.300 ;
        RECT 30.940 48.000 31.900 57.190 ;
        RECT 34.720 57.170 35.800 57.190 ;
        RECT 38.870 57.170 39.950 57.190 ;
        RECT 40.880 56.340 41.840 57.190 ;
        RECT 44.660 57.150 45.620 57.210 ;
        RECT 32.860 54.030 33.820 56.300 ;
        RECT 27.595 47.670 30.620 48.000 ;
        RECT 27.645 47.640 27.975 47.670 ;
        RECT 6.260 45.390 24.910 46.590 ;
        RECT 6.170 35.170 7.490 36.370 ;
        RECT 23.710 35.180 24.910 45.390 ;
        RECT 30.290 44.400 30.620 47.670 ;
        RECT 30.930 44.400 31.900 48.000 ;
        RECT 30.300 43.890 30.620 44.400 ;
        RECT 30.940 43.890 31.900 44.400 ;
        RECT 30.290 43.290 30.620 43.890 ;
        RECT 30.290 40.290 30.610 43.290 ;
        RECT 30.930 42.020 31.900 43.890 ;
        RECT 32.850 52.700 33.820 54.030 ;
        RECT 32.850 52.190 33.810 52.700 ;
        RECT 32.850 48.590 33.820 52.190 ;
        RECT 37.645 48.715 38.035 49.045 ;
        RECT 30.930 40.290 31.890 42.020 ;
        RECT 32.850 38.110 33.810 48.590 ;
        RECT 37.675 48.040 38.005 48.715 ;
        RECT 40.210 48.040 40.530 56.340 ;
        RECT 40.850 55.000 41.840 56.340 ;
        RECT 40.850 53.800 41.810 55.000 ;
        RECT 37.505 47.710 40.530 48.040 ;
        RECT 40.200 44.440 40.530 47.710 ;
        RECT 40.210 43.930 40.530 44.440 ;
        RECT 40.200 43.460 40.530 43.930 ;
        RECT 40.840 52.740 41.810 53.800 ;
        RECT 40.840 52.230 41.800 52.740 ;
        RECT 40.840 48.630 41.810 52.230 ;
        RECT 40.200 40.330 40.520 43.460 ;
        RECT 40.840 40.330 41.800 48.630 ;
        RECT 42.770 48.040 43.730 56.340 ;
        RECT 42.760 44.440 43.730 48.040 ;
        RECT 46.440 45.220 53.770 59.290 ;
        RECT 55.830 52.890 56.150 58.060 ;
        RECT 56.470 54.460 57.430 59.290 ;
        RECT 60.280 59.270 61.240 59.290 ;
        RECT 58.390 51.410 59.350 58.060 ;
        RECT 64.300 57.900 64.660 61.500 ;
        RECT 64.970 57.900 65.940 61.500 ;
        RECT 66.890 57.900 67.860 61.500 ;
        RECT 75.470 58.460 75.790 63.440 ;
        RECT 76.100 62.880 77.060 63.440 ;
        RECT 76.100 60.630 77.070 62.880 ;
        RECT 76.110 59.280 77.070 60.630 ;
        RECT 78.030 58.660 78.990 63.440 ;
        RECT 84.820 58.660 85.140 62.880 ;
        RECT 85.460 59.280 86.420 65.370 ;
        RECT 89.300 65.020 90.260 65.370 ;
        RECT 89.240 64.060 90.320 65.020 ;
        RECT 78.030 58.460 85.140 58.660 ;
        RECT 75.470 58.140 85.140 58.460 ;
        RECT 64.300 57.370 64.620 57.900 ;
        RECT 64.300 54.230 64.650 57.370 ;
        RECT 64.330 51.410 64.650 54.230 ;
        RECT 64.970 52.610 65.930 57.900 ;
        RECT 64.940 51.650 65.960 52.610 ;
        RECT 66.890 51.520 67.850 57.900 ;
        RECT 78.030 57.700 85.140 58.140 ;
        RECT 78.030 57.360 78.990 57.700 ;
        RECT 75.400 51.520 75.720 57.360 ;
        RECT 76.040 52.220 77.000 57.360 ;
        RECT 77.960 55.350 78.990 57.360 ;
        RECT 87.380 55.525 88.340 62.880 ;
        RECT 104.125 55.525 104.455 55.555 ;
        RECT 77.960 53.760 78.920 55.350 ;
        RECT 87.315 55.195 104.455 55.525 ;
        RECT 87.380 54.620 88.340 55.195 ;
        RECT 104.125 55.165 104.455 55.195 ;
        RECT 108.740 55.250 109.940 66.690 ;
        RECT 126.290 66.660 127.490 66.720 ;
        RECT 137.410 64.830 137.730 66.720 ;
        RECT 138.050 64.830 139.010 66.360 ;
        RECT 139.970 64.830 140.930 66.720 ;
        RECT 137.400 64.090 137.730 64.830 ;
        RECT 137.400 61.700 137.720 64.090 ;
        RECT 138.040 63.160 139.010 64.830 ;
        RECT 139.960 63.520 140.930 64.830 ;
        RECT 138.040 62.150 139.000 63.160 ;
        RECT 137.400 61.230 137.750 61.700 ;
        RECT 138.040 61.230 139.030 62.150 ;
        RECT 139.960 61.230 140.920 63.520 ;
        RECT 137.430 59.810 137.750 61.230 ;
        RECT 138.070 59.810 139.030 61.230 ;
        RECT 137.420 58.580 137.750 59.810 ;
        RECT 137.420 56.210 137.740 58.580 ;
        RECT 138.060 57.700 139.030 59.810 ;
        RECT 138.060 56.210 139.020 57.700 ;
        RECT 139.980 56.670 140.940 59.810 ;
        RECT 139.980 56.210 140.950 56.670 ;
        RECT 108.740 54.050 127.300 55.250 ;
        RECT 90.210 52.980 92.430 53.330 ;
        RECT 90.210 52.660 97.200 52.980 ;
        RECT 90.210 52.110 92.430 52.660 ;
        RECT 66.890 51.410 75.840 51.520 ;
        RECT 58.390 50.560 75.840 51.410 ;
        RECT 58.390 50.480 67.850 50.560 ;
        RECT 58.430 50.450 67.850 50.480 ;
        RECT 71.790 49.120 72.990 49.180 ;
        RECT 64.060 48.455 72.990 49.120 ;
        RECT 62.900 48.125 72.990 48.455 ;
        RECT 64.040 47.920 72.990 48.125 ;
        RECT 60.200 45.220 61.160 45.230 ;
        RECT 46.440 44.670 63.090 45.220 ;
        RECT 42.770 43.930 43.730 44.440 ;
        RECT 46.560 44.260 63.090 44.670 ;
        RECT 42.760 42.400 43.730 43.930 ;
        RECT 52.470 42.780 53.430 44.260 ;
        RECT 60.200 44.020 61.160 44.260 ;
        RECT 62.120 44.220 63.090 44.260 ;
        RECT 60.140 43.060 61.220 44.020 ;
        RECT 42.760 38.460 43.720 42.400 ;
        RECT 61.480 39.310 61.800 42.450 ;
        RECT 62.120 40.600 63.080 44.220 ;
        RECT 61.480 38.850 61.810 39.310 ;
        RECT 62.120 38.850 63.090 40.600 ;
        RECT 64.040 38.850 65.000 47.920 ;
        RECT 71.790 47.860 72.990 47.920 ;
        RECT 77.720 49.120 78.920 49.180 ;
        RECT 77.720 49.110 80.560 49.120 ;
        RECT 81.510 49.110 82.710 49.170 ;
        RECT 77.720 47.910 82.710 49.110 ;
        RECT 77.720 47.860 78.920 47.910 ;
        RECT 81.510 47.850 82.710 47.910 ;
        RECT 30.300 38.060 33.890 38.110 ;
        RECT 30.300 37.790 40.540 38.060 ;
        RECT 6.230 19.400 7.430 35.170 ;
        RECT 30.300 32.530 30.620 37.790 ;
        RECT 32.850 37.740 40.540 37.790 ;
        RECT 32.850 36.130 33.810 37.740 ;
        RECT 30.940 30.430 31.900 36.130 ;
        RECT 32.850 34.130 33.820 36.130 ;
        RECT 32.860 32.530 33.820 34.130 ;
        RECT 40.220 32.520 40.540 37.740 ;
        RECT 42.760 37.500 57.210 38.460 ;
        RECT 42.760 36.120 43.720 37.500 ;
        RECT 40.860 30.550 41.820 36.120 ;
        RECT 42.760 34.250 43.740 36.120 ;
        RECT 42.780 32.520 43.740 34.250 ;
        RECT 56.890 34.420 57.210 37.500 ;
        RECT 61.490 34.420 61.810 38.850 ;
        RECT 62.130 34.730 63.090 38.850 ;
        RECT 56.890 34.100 61.810 34.420 ;
        RECT 61.490 32.570 61.810 34.100 ;
        RECT 50.115 24.040 53.165 24.225 ;
        RECT 64.050 24.040 65.010 38.330 ;
        RECT 87.410 30.950 88.610 30.960 ;
        RECT 50.115 23.080 65.010 24.040 ;
        RECT 50.115 21.175 53.165 23.080 ;
        RECT 64.050 22.750 65.010 23.080 ;
        RECT 66.730 30.940 90.390 30.950 ;
        RECT 91.680 30.940 92.880 49.100 ;
        RECT 66.730 20.800 92.880 30.940 ;
        RECT 96.880 22.350 97.200 52.660 ;
        RECT 108.610 43.050 109.810 50.390 ;
        RECT 126.100 49.100 127.300 54.050 ;
        RECT 131.310 54.610 134.820 54.660 ;
        RECT 139.990 54.610 140.950 56.210 ;
        RECT 147.010 54.630 147.970 54.690 ;
        RECT 142.490 54.610 147.970 54.630 ;
        RECT 131.310 53.700 147.970 54.610 ;
        RECT 133.290 53.670 147.970 53.700 ;
        RECT 133.290 53.650 144.190 53.670 ;
        RECT 129.995 44.460 130.325 45.515 ;
        RECT 132.650 44.460 132.970 52.760 ;
        RECT 133.290 44.460 134.250 53.650 ;
        RECT 137.070 53.630 138.150 53.650 ;
        RECT 141.220 53.630 142.300 53.650 ;
        RECT 143.230 52.800 144.190 53.650 ;
        RECT 147.010 53.610 147.970 53.670 ;
        RECT 135.210 50.490 136.170 52.760 ;
        RECT 129.945 44.130 132.970 44.460 ;
        RECT 108.610 41.850 127.260 43.050 ;
        RECT 108.520 31.630 109.840 32.830 ;
        RECT 126.060 31.640 127.260 41.850 ;
        RECT 132.640 40.860 132.970 44.130 ;
        RECT 133.280 40.860 134.250 44.460 ;
        RECT 132.650 40.350 132.970 40.860 ;
        RECT 133.290 40.350 134.250 40.860 ;
        RECT 132.640 39.750 132.970 40.350 ;
        RECT 132.640 36.750 132.960 39.750 ;
        RECT 133.280 38.480 134.250 40.350 ;
        RECT 135.200 49.160 136.170 50.490 ;
        RECT 135.200 48.650 136.160 49.160 ;
        RECT 135.200 45.050 136.170 48.650 ;
        RECT 133.280 36.750 134.240 38.480 ;
        RECT 135.200 34.570 136.160 45.050 ;
        RECT 139.865 44.500 140.195 44.530 ;
        RECT 142.560 44.500 142.880 52.800 ;
        RECT 143.200 51.460 144.190 52.800 ;
        RECT 143.200 50.260 144.160 51.460 ;
        RECT 139.855 44.170 142.880 44.500 ;
        RECT 139.865 44.140 140.195 44.170 ;
        RECT 142.550 40.900 142.880 44.170 ;
        RECT 142.560 40.390 142.880 40.900 ;
        RECT 142.550 39.920 142.880 40.390 ;
        RECT 143.190 49.200 144.160 50.260 ;
        RECT 143.190 48.690 144.150 49.200 ;
        RECT 143.190 45.090 144.160 48.690 ;
        RECT 142.550 36.790 142.870 39.920 ;
        RECT 143.190 36.790 144.150 45.090 ;
        RECT 145.120 44.500 146.080 52.800 ;
        RECT 145.110 40.900 146.080 44.500 ;
        RECT 145.120 40.390 146.080 40.900 ;
        RECT 145.110 38.860 146.080 40.390 ;
        RECT 145.110 34.920 146.070 38.860 ;
        RECT 150.830 34.920 151.790 37.230 ;
        RECT 132.650 34.520 136.240 34.570 ;
        RECT 132.650 34.250 142.890 34.520 ;
        RECT 97.520 22.350 98.480 25.950 ;
        RECT 98.800 22.350 99.760 28.590 ;
        RECT 88.390 20.720 92.880 20.800 ;
        RECT 91.680 20.700 92.880 20.720 ;
        RECT 97.640 20.540 98.480 22.350 ;
        RECT 103.040 19.950 104.360 22.010 ;
        RECT 4.520 18.850 5.080 18.910 ;
        RECT 6.230 18.850 30.090 19.400 ;
        RECT 4.520 18.290 30.090 18.850 ;
        RECT 102.980 18.630 104.420 19.950 ;
        RECT 4.520 18.230 5.080 18.290 ;
        RECT 6.230 18.200 30.090 18.290 ;
        RECT 108.580 15.860 109.780 31.630 ;
        RECT 132.650 28.990 132.970 34.250 ;
        RECT 135.200 34.200 142.890 34.250 ;
        RECT 135.200 32.590 136.160 34.200 ;
        RECT 133.290 26.890 134.250 32.590 ;
        RECT 135.200 30.590 136.170 32.590 ;
        RECT 135.210 28.990 136.170 30.590 ;
        RECT 142.570 28.980 142.890 34.200 ;
        RECT 145.110 33.960 159.290 34.920 ;
        RECT 145.110 32.580 146.070 33.960 ;
        RECT 143.210 27.010 144.170 32.580 ;
        RECT 145.110 30.710 146.090 32.580 ;
        RECT 145.130 28.980 146.090 30.710 ;
        RECT 106.870 15.310 107.430 15.370 ;
        RECT 108.580 15.310 132.440 15.860 ;
        RECT 106.870 14.750 132.440 15.310 ;
        RECT 106.870 14.690 107.430 14.750 ;
        RECT 108.580 14.660 132.440 14.750 ;
      LAYER met2 ;
        RECT 59.300 204.370 60.260 204.400 ;
        RECT 59.300 203.410 64.145 204.370 ;
        RECT 59.300 203.380 60.260 203.410 ;
        RECT 53.495 195.910 60.290 196.870 ;
        RECT 53.420 188.790 60.620 189.990 ;
        RECT 63.620 189.600 108.120 190.290 ;
        RECT 63.620 189.090 108.130 189.600 ;
        RECT 38.740 186.550 39.060 188.595 ;
        RECT 53.420 186.550 54.620 188.790 ;
        RECT 38.710 186.230 39.090 186.550 ;
        RECT 47.710 186.230 54.620 186.550 ;
        RECT 53.420 164.790 54.620 186.230 ;
        RECT 63.620 186.550 64.820 189.090 ;
        RECT 78.980 186.550 79.300 188.595 ;
        RECT 63.620 186.230 70.330 186.550 ;
        RECT 78.950 186.230 79.330 186.550 ;
        RECT 63.620 185.890 64.820 186.230 ;
        RECT 106.920 176.200 108.130 189.090 ;
        RECT 106.920 175.190 117.650 176.200 ;
        RECT 107.110 175.180 117.650 175.190 ;
        RECT 55.860 166.550 56.180 166.580 ;
        RECT 55.860 166.230 57.225 166.550 ;
        RECT 55.860 166.200 56.180 166.230 ;
        RECT 36.170 164.490 63.170 164.790 ;
        RECT 35.920 160.250 37.120 160.280 ;
        RECT 35.920 159.050 43.965 160.250 ;
        RECT 35.920 159.020 37.120 159.050 ;
        RECT 52.680 158.440 52.960 158.475 ;
        RECT 51.140 158.140 52.970 158.440 ;
        RECT 52.680 158.105 52.960 158.140 ;
        RECT 53.420 150.990 54.620 164.490 ;
        RECT 64.840 159.670 65.800 159.700 ;
        RECT 64.840 158.710 67.645 159.670 ;
        RECT 64.840 158.680 65.800 158.710 ;
        RECT 66.740 157.440 67.620 157.780 ;
        RECT 69.440 157.440 70.320 157.780 ;
        RECT 65.910 156.040 66.270 156.340 ;
        RECT 69.440 156.305 71.990 156.330 ;
        RECT 65.940 154.540 66.240 156.040 ;
        RECT 69.420 155.475 71.990 156.305 ;
        RECT 69.440 155.450 71.990 155.475 ;
        RECT 65.940 154.240 72.170 154.540 ;
        RECT 65.370 154.040 65.670 154.070 ;
        RECT 61.370 153.930 65.670 154.040 ;
        RECT 48.890 149.790 54.620 150.990 ;
        RECT 61.240 153.740 65.670 153.930 ;
        RECT 61.240 133.190 61.560 153.740 ;
        RECT 65.370 153.710 65.670 153.740 ;
        RECT 65.920 152.340 66.800 152.680 ;
        RECT 68.620 152.340 69.500 152.680 ;
        RECT 64.120 151.440 65.000 151.480 ;
        RECT 64.120 151.140 65.620 151.440 ;
        RECT 65.320 148.240 65.620 151.140 ;
        RECT 68.620 149.940 69.500 150.280 ;
        RECT 65.920 149.140 66.800 149.480 ;
        RECT 70.420 148.240 71.300 148.280 ;
        RECT 65.320 147.940 71.300 148.240 ;
        RECT 65.920 146.740 66.800 147.080 ;
        RECT 68.620 146.740 69.500 147.080 ;
        RECT 65.920 145.140 66.800 145.480 ;
        RECT 68.620 145.140 69.500 145.480 ;
        RECT 65.920 142.740 66.800 143.080 ;
        RECT 68.620 142.740 69.500 143.080 ;
        RECT 65.920 140.340 66.800 140.680 ;
        RECT 68.620 140.340 69.500 140.680 ;
        RECT 71.870 140.040 72.170 154.240 ;
        RECT 100.920 152.490 102.120 152.520 ;
        RECT 98.875 151.290 102.120 152.490 ;
        RECT 100.920 151.260 102.120 151.290 ;
        RECT 70.840 139.740 72.170 140.040 ;
        RECT 65.920 138.740 66.800 139.080 ;
        RECT 68.620 138.740 69.500 139.080 ;
        RECT 68.620 137.940 69.500 138.280 ;
        RECT 65.920 136.340 66.800 136.680 ;
        RECT 68.620 136.340 69.500 136.680 ;
        RECT 65.920 135.540 66.800 135.880 ;
        RECT 68.620 135.540 69.500 135.880 ;
        RECT 65.920 134.740 66.800 135.080 ;
        RECT 68.620 134.740 69.500 135.080 ;
        RECT 61.170 132.740 61.620 133.190 ;
        RECT 66.440 133.130 67.400 133.160 ;
        RECT 66.440 132.170 70.345 133.130 ;
        RECT 66.440 132.140 67.400 132.170 ;
        RECT 66.730 131.815 67.610 131.840 ;
        RECT 66.710 130.985 67.630 131.815 ;
        RECT 66.730 129.110 67.610 130.985 ;
        RECT 104.095 55.195 104.485 55.525 ;
        RECT 58.650 53.240 58.970 53.245 ;
        RECT 55.800 52.920 58.970 53.240 ;
        RECT 58.650 52.875 58.970 52.920 ;
        RECT 27.645 51.165 63.260 51.495 ;
        RECT 27.645 48.000 27.975 51.165 ;
        RECT 37.675 50.225 58.655 50.555 ;
        RECT 37.675 48.685 38.005 50.225 ;
        RECT 27.615 47.670 28.005 48.000 ;
        RECT 52.440 42.810 53.460 43.770 ;
        RECT 52.470 41.155 53.430 42.810 ;
        RECT 58.325 33.795 58.655 50.225 ;
        RECT 62.930 48.095 63.260 51.165 ;
        RECT 104.125 45.485 104.455 55.195 ;
        RECT 111.005 49.715 111.335 81.335 ;
        RECT 111.005 49.385 140.195 49.715 ;
        RECT 101.960 45.155 130.355 45.485 ;
        RECT 139.865 44.500 140.195 49.385 ;
        RECT 139.835 44.170 140.225 44.500 ;
        RECT 58.325 33.465 64.765 33.795 ;
        RECT 59.925 32.600 61.840 32.920 ;
        RECT 98.800 28.560 99.760 30.645 ;
        RECT 98.770 27.600 99.790 28.560 ;
        RECT 103.040 21.980 104.360 23.965 ;
        RECT 103.010 20.660 104.390 21.980 ;
      LAYER met3 ;
        RECT 38.715 188.570 39.085 188.575 ;
        RECT 53.420 188.570 54.620 196.990 ;
        RECT 38.715 188.250 54.620 188.570 ;
        RECT 38.715 188.245 39.085 188.250 ;
        RECT 42.745 160.250 43.945 160.275 ;
        RECT 53.420 160.250 54.620 188.250 ;
        RECT 63.165 188.970 64.125 204.395 ;
        RECT 63.165 188.010 82.700 188.970 ;
        RECT 56.875 166.550 57.205 166.575 ;
        RECT 56.860 166.230 59.680 166.550 ;
        RECT 56.875 166.205 57.205 166.230 ;
        RECT 59.360 164.790 59.680 166.230 ;
        RECT 42.745 159.050 54.620 160.250 ;
        RECT 56.120 159.390 61.520 164.790 ;
        RECT 42.745 159.025 43.945 159.050 ;
        RECT 52.655 158.440 52.985 158.455 ;
        RECT 54.960 158.440 55.280 158.480 ;
        RECT 52.655 158.140 55.280 158.440 ;
        RECT 52.655 158.125 52.985 158.140 ;
        RECT 54.960 158.100 55.280 158.140 ;
        RECT 66.665 155.270 67.625 159.695 ;
        RECT 69.440 155.450 70.320 158.790 ;
        RECT 66.665 154.830 69.200 155.270 ;
        RECT 66.665 154.310 69.500 154.830 ;
        RECT 65.920 131.840 66.800 153.690 ;
        RECT 68.620 134.490 69.500 154.310 ;
        RECT 81.740 151.590 82.700 188.010 ;
        RECT 98.895 152.490 100.095 152.515 ;
        RECT 79.020 146.190 84.420 151.590 ;
        RECT 86.820 146.190 92.220 151.590 ;
        RECT 96.890 151.290 100.095 152.490 ;
        RECT 98.895 151.265 100.095 151.290 ;
        RECT 81.520 143.790 81.920 146.190 ;
        RECT 89.320 143.790 89.720 146.190 ;
        RECT 79.020 140.370 84.420 143.790 ;
        RECT 74.540 139.410 84.420 140.370 ;
        RECT 69.365 133.130 70.325 133.155 ;
        RECT 74.540 133.130 75.500 139.410 ;
        RECT 79.020 138.890 84.420 139.410 ;
        RECT 86.820 138.890 92.220 143.790 ;
        RECT 79.020 138.390 92.220 138.890 ;
        RECT 69.365 132.170 75.500 133.130 ;
        RECT 69.365 132.145 70.325 132.170 ;
        RECT 65.920 130.960 67.610 131.840 ;
        RECT 58.625 52.895 58.995 53.225 ;
        RECT 52.445 41.175 53.455 42.135 ;
        RECT 52.470 36.720 53.430 41.175 ;
        RECT 50.560 31.320 55.960 36.720 ;
        RECT 58.650 32.920 58.970 52.895 ;
        RECT 101.980 45.485 102.310 45.510 ;
        RECT 100.485 45.130 102.310 45.485 ;
        RECT 100.485 42.310 100.815 45.130 ;
        RECT 98.080 36.910 103.480 42.310 ;
        RECT 59.945 32.920 60.275 32.945 ;
        RECT 58.270 32.600 60.275 32.920 ;
        RECT 58.650 32.570 58.970 32.600 ;
        RECT 59.945 32.575 60.275 32.600 ;
        RECT 98.800 30.625 99.760 36.910 ;
        RECT 98.775 29.665 99.785 30.625 ;
        RECT 103.040 23.945 104.360 26.250 ;
        RECT 103.015 22.625 104.385 23.945 ;
      LAYER met4 ;
        RECT 56.120 159.390 61.520 164.790 ;
        RECT 54.955 158.440 55.285 158.455 ;
        RECT 57.570 158.440 57.870 159.390 ;
        RECT 54.955 158.140 57.870 158.440 ;
        RECT 54.955 158.125 55.285 158.140 ;
        RECT 79.020 146.190 84.420 151.590 ;
        RECT 86.820 150.490 92.220 151.590 ;
        RECT 96.915 150.490 98.115 152.495 ;
        RECT 86.820 149.290 98.115 150.490 ;
        RECT 86.820 146.190 92.220 149.290 ;
        RECT 81.520 143.790 81.920 146.190 ;
        RECT 89.320 143.790 89.720 146.190 ;
        RECT 79.020 138.890 84.420 143.790 ;
        RECT 86.820 138.890 92.220 143.790 ;
        RECT 79.020 138.390 92.220 138.890 ;
        RECT 98.080 42.280 103.480 42.310 ;
        RECT 98.080 36.910 104.360 42.280 ;
        RECT 50.560 32.920 55.960 36.720 ;
        RECT 58.295 32.920 58.625 32.925 ;
        RECT 50.560 32.600 58.625 32.920 ;
        RECT 50.560 31.320 55.960 32.600 ;
        RECT 58.295 32.595 58.625 32.600 ;
        RECT 103.040 26.225 104.360 36.910 ;
        RECT 103.035 24.905 104.365 26.225 ;
  END
END tt_um_jnw_wulffern
END LIBRARY

