MACRO tt_um_jnw_wulffern
  CLASS BLOCK ;
  FOREIGN tt_um_jnw_wulffern ;
  ORIGIN -0.580 -5.000 ;
  SIZE 161.680 BY 220.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.288000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.288000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.936000 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.936000 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.044000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 51.500 204.790 59.100 210.070 ;
        RECT 60.500 204.290 68.100 209.570 ;
        RECT 69.500 204.290 77.100 209.570 ;
        RECT 78.500 204.290 86.100 209.570 ;
        RECT 96.500 204.290 104.100 209.570 ;
        RECT 114.900 204.290 122.500 209.570 ;
        RECT 123.900 204.290 131.500 209.570 ;
        RECT 132.900 204.290 140.500 209.570 ;
        RECT 141.900 204.790 149.500 210.070 ;
        RECT 51.500 197.290 59.100 202.570 ;
        RECT 60.500 197.290 68.100 202.570 ;
        RECT 69.500 197.290 77.100 202.570 ;
        RECT 78.500 197.290 86.100 202.570 ;
        RECT 87.500 197.290 95.100 202.570 ;
        RECT 96.500 197.290 104.100 202.570 ;
        RECT 105.900 197.290 113.500 202.570 ;
        RECT 114.900 197.290 122.500 202.570 ;
        RECT 123.900 197.290 131.500 202.570 ;
        RECT 132.900 197.290 140.500 202.570 ;
        RECT 141.900 197.290 149.500 202.570 ;
      LAYER pwell ;
        RECT 152.320 195.690 158.080 210.090 ;
      LAYER nwell ;
        RECT 51.500 190.290 59.100 195.570 ;
        RECT 60.500 190.290 68.100 195.570 ;
        RECT 69.500 190.290 77.100 195.570 ;
        RECT 78.500 190.290 86.100 195.570 ;
        RECT 96.500 190.290 104.100 195.570 ;
        RECT 114.900 190.290 122.500 195.570 ;
        RECT 123.900 190.290 131.500 195.570 ;
        RECT 132.900 190.290 140.500 195.570 ;
        RECT 141.900 190.290 149.500 195.570 ;
      LAYER pwell ;
        RECT 56.320 172.690 75.040 187.090 ;
      LAYER nwell ;
        RECT 78.500 181.790 86.100 187.070 ;
        RECT 87.500 181.290 95.100 186.570 ;
        RECT 105.900 181.290 113.500 186.570 ;
        RECT 114.900 181.790 122.500 187.070 ;
        RECT 78.500 174.290 86.100 179.570 ;
        RECT 87.500 174.290 95.100 179.570 ;
        RECT 105.900 174.290 113.500 179.570 ;
        RECT 114.900 174.290 122.500 179.570 ;
      LAYER pwell ;
        RECT 125.960 172.690 144.680 187.090 ;
        RECT 152.320 177.690 158.080 192.090 ;
        RECT 16.690 149.630 22.390 167.630 ;
      LAYER nwell ;
        RECT 22.390 149.630 28.090 167.630 ;
      LAYER pwell ;
        RECT 56.320 154.690 75.040 169.090 ;
        RECT 78.500 161.290 86.100 171.570 ;
        RECT 87.500 161.290 95.100 171.570 ;
        RECT 105.900 161.290 113.500 171.570 ;
        RECT 114.900 161.290 122.500 171.570 ;
        RECT 79.500 157.225 86.200 157.990 ;
        RECT 79.500 152.055 80.265 157.225 ;
        RECT 85.435 152.055 86.200 157.225 ;
        RECT 79.500 151.290 86.200 152.055 ;
        RECT 87.500 157.225 94.200 157.990 ;
        RECT 87.500 152.055 88.265 157.225 ;
        RECT 93.435 152.055 94.200 157.225 ;
        RECT 87.500 151.290 94.200 152.055 ;
        RECT 95.500 157.225 102.200 157.990 ;
        RECT 95.500 152.055 96.265 157.225 ;
        RECT 101.435 152.055 102.200 157.225 ;
      LAYER nwell ;
        RECT 104.300 155.690 110.000 159.290 ;
      LAYER pwell ;
        RECT 110.000 155.690 115.700 159.290 ;
        RECT 125.960 154.690 144.680 169.090 ;
        RECT 152.320 159.690 158.080 174.090 ;
        RECT 95.500 151.290 102.200 152.055 ;
        RECT 56.320 136.690 75.040 151.090 ;
        RECT 79.500 149.225 86.200 149.990 ;
        RECT 79.500 144.055 80.265 149.225 ;
        RECT 85.435 144.055 86.200 149.225 ;
        RECT 79.500 143.290 86.200 144.055 ;
        RECT 87.500 149.225 94.200 149.990 ;
        RECT 87.500 144.055 88.265 149.225 ;
        RECT 93.435 144.055 94.200 149.225 ;
        RECT 87.500 143.290 94.200 144.055 ;
        RECT 95.500 149.225 102.200 149.990 ;
        RECT 95.500 144.055 96.265 149.225 ;
        RECT 101.435 144.055 102.200 149.225 ;
        RECT 95.500 143.290 102.200 144.055 ;
        RECT 79.500 141.225 86.200 141.990 ;
        RECT 79.500 136.055 80.265 141.225 ;
        RECT 85.435 136.055 86.200 141.225 ;
        RECT 79.500 135.290 86.200 136.055 ;
        RECT 87.500 141.225 94.200 141.990 ;
        RECT 87.500 136.055 88.265 141.225 ;
        RECT 93.435 136.055 94.200 141.225 ;
        RECT 87.500 135.290 94.200 136.055 ;
        RECT 95.500 141.225 102.200 141.990 ;
        RECT 95.500 136.055 96.265 141.225 ;
        RECT 101.435 136.055 102.200 141.225 ;
        RECT 95.500 135.290 102.200 136.055 ;
        RECT 103.500 133.870 109.200 154.190 ;
        RECT 101.000 133.790 109.200 133.870 ;
      LAYER nwell ;
        RECT 109.200 133.790 114.900 154.190 ;
      LAYER pwell ;
        RECT 152.320 141.690 158.080 156.090 ;
        RECT 56.320 118.690 75.040 133.090 ;
        RECT 80.320 118.690 99.040 133.090 ;
        RECT 101.000 123.790 107.960 133.790 ;
      LAYER nwell ;
        RECT 73.850 97.380 81.450 101.540 ;
        RECT 73.830 96.260 81.450 97.380 ;
      LAYER pwell ;
        RECT 62.690 91.490 70.290 95.620 ;
      LAYER nwell ;
        RECT 73.830 93.390 81.430 96.260 ;
        RECT 73.830 92.100 81.470 93.390 ;
      LAYER pwell ;
        RECT 62.680 90.340 70.290 91.490 ;
        RECT 62.680 87.490 70.280 90.340 ;
      LAYER nwell ;
        RECT 73.870 89.230 81.470 92.100 ;
        RECT 73.830 88.110 81.470 89.230 ;
      LAYER pwell ;
        RECT 62.680 86.210 70.310 87.490 ;
        RECT 62.710 83.360 70.310 86.210 ;
      LAYER nwell ;
        RECT 73.830 85.230 81.430 88.110 ;
      LAYER pwell ;
        RECT 92.410 86.600 98.170 101.000 ;
        RECT 103.080 86.680 108.840 101.080 ;
        RECT 113.670 86.760 119.430 101.160 ;
      LAYER nwell ;
        RECT 73.830 83.950 81.450 85.230 ;
      LAYER pwell ;
        RECT 62.700 82.210 70.310 83.360 ;
        RECT 62.700 79.370 70.300 82.210 ;
      LAYER nwell ;
        RECT 73.850 81.070 81.450 83.950 ;
        RECT 73.830 79.950 81.450 81.070 ;
      LAYER pwell ;
        RECT 62.700 78.080 70.310 79.370 ;
        RECT 62.710 75.240 70.310 78.080 ;
      LAYER nwell ;
        RECT 73.830 76.940 81.430 79.950 ;
        RECT 73.830 75.790 81.450 76.940 ;
      LAYER pwell ;
        RECT 62.700 74.090 70.310 75.240 ;
        RECT 6.500 57.830 25.220 72.230 ;
        RECT 62.700 71.230 70.300 74.090 ;
      LAYER nwell ;
        RECT 73.850 72.780 81.450 75.790 ;
        RECT 73.850 71.660 81.460 72.780 ;
        RECT 33.440 64.960 41.040 69.980 ;
      LAYER pwell ;
        RECT 62.700 69.960 70.330 71.230 ;
        RECT 62.730 67.100 70.330 69.960 ;
      LAYER nwell ;
        RECT 73.860 68.650 81.460 71.660 ;
      LAYER pwell ;
        RECT 62.720 65.950 70.330 67.100 ;
      LAYER nwell ;
        RECT 73.840 67.500 81.460 68.650 ;
        RECT 33.440 64.700 41.060 64.960 ;
        RECT 33.460 59.680 41.060 64.700 ;
      LAYER pwell ;
        RECT 62.720 63.110 70.320 65.950 ;
      LAYER nwell ;
        RECT 73.840 64.490 81.440 67.500 ;
        RECT 73.840 63.370 81.460 64.490 ;
      LAYER pwell ;
        RECT 62.720 61.820 70.330 63.110 ;
        RECT 6.400 40.240 25.120 54.640 ;
      LAYER nwell ;
        RECT 28.690 49.610 36.290 57.910 ;
        RECT 38.600 49.650 46.200 57.950 ;
        RECT 54.220 54.390 61.820 59.670 ;
      LAYER pwell ;
        RECT 62.730 58.980 70.330 61.820 ;
      LAYER nwell ;
        RECT 73.860 59.210 81.460 63.370 ;
        RECT 83.210 59.210 90.810 64.490 ;
      LAYER pwell ;
        RECT 62.720 57.830 70.330 58.980 ;
        RECT 62.720 53.700 70.320 57.830 ;
        RECT 73.790 53.690 81.390 58.970 ;
        RECT 108.850 54.290 127.570 68.690 ;
      LAYER nwell ;
        RECT 135.790 61.420 143.390 66.440 ;
        RECT 135.790 61.160 143.410 61.420 ;
        RECT 135.810 56.140 143.410 61.160 ;
        RECT 28.680 48.520 36.290 49.610 ;
        RECT 38.590 48.560 46.200 49.650 ;
        RECT 28.680 40.220 36.280 48.520 ;
        RECT 38.590 40.260 46.190 48.560 ;
        RECT 59.870 39.940 67.470 44.060 ;
        RECT 59.870 38.780 67.480 39.940 ;
      LAYER pwell ;
        RECT 6.340 22.770 25.060 37.170 ;
        RECT 28.690 32.460 36.290 37.740 ;
        RECT 38.610 32.450 46.210 37.730 ;
      LAYER nwell ;
        RECT 59.880 34.660 67.480 38.780 ;
      LAYER pwell ;
        RECT 72.600 35.490 78.360 49.890 ;
        RECT 82.370 35.410 92.450 49.810 ;
        RECT 108.750 36.700 127.470 51.100 ;
      LAYER nwell ;
        RECT 131.040 46.070 138.640 54.370 ;
        RECT 140.950 46.110 148.550 54.410 ;
        RECT 131.030 44.980 138.640 46.070 ;
        RECT 140.940 45.020 148.550 46.110 ;
        RECT 131.030 36.680 138.630 44.980 ;
        RECT 140.940 36.720 148.540 45.020 ;
      LAYER pwell ;
        RECT 68.170 29.815 74.870 30.580 ;
        RECT 68.170 24.645 68.935 29.815 ;
        RECT 74.105 24.645 74.870 29.815 ;
        RECT 68.170 23.880 74.870 24.645 ;
        RECT 76.140 29.815 82.840 30.580 ;
        RECT 76.140 24.645 76.905 29.815 ;
        RECT 82.075 24.645 82.840 29.815 ;
        RECT 76.140 23.880 82.840 24.645 ;
        RECT 84.110 29.815 90.810 30.580 ;
        RECT 84.110 24.645 84.875 29.815 ;
        RECT 90.045 24.645 90.810 29.815 ;
        RECT 84.110 23.880 90.810 24.645 ;
        RECT 68.170 21.715 74.870 22.480 ;
        RECT 68.170 16.545 68.935 21.715 ;
        RECT 74.105 16.545 74.870 21.715 ;
        RECT 68.170 15.780 74.870 16.545 ;
        RECT 76.140 21.715 82.840 22.480 ;
        RECT 76.140 16.545 76.905 21.715 ;
        RECT 82.075 16.545 82.840 21.715 ;
        RECT 76.140 15.780 82.840 16.545 ;
        RECT 84.110 21.715 90.810 22.480 ;
        RECT 95.270 22.280 102.230 27.560 ;
        RECT 84.110 16.545 84.875 21.715 ;
        RECT 90.045 16.545 90.810 21.715 ;
        RECT 108.690 19.230 127.410 33.630 ;
        RECT 131.040 28.920 138.640 34.200 ;
        RECT 140.960 28.910 148.560 34.190 ;
        RECT 84.110 15.780 90.810 16.545 ;
        RECT 68.170 13.615 74.870 14.380 ;
        RECT 68.170 8.445 68.935 13.615 ;
        RECT 74.105 8.445 74.870 13.615 ;
        RECT 68.170 7.680 74.870 8.445 ;
        RECT 76.140 13.615 82.840 14.380 ;
        RECT 76.140 8.445 76.905 13.615 ;
        RECT 82.075 8.445 82.840 13.615 ;
        RECT 76.140 7.680 82.840 8.445 ;
        RECT 84.110 13.615 90.810 14.380 ;
        RECT 84.110 8.445 84.875 13.615 ;
        RECT 90.045 8.445 90.810 13.615 ;
        RECT 84.110 7.680 90.810 8.445 ;
      LAYER li1 ;
        RECT 52.000 210.770 149.000 211.790 ;
        RECT 150.500 210.850 160.500 211.790 ;
        RECT 51.940 209.810 149.060 210.770 ;
        RECT 51.940 190.770 52.900 209.810 ;
        RECT 53.860 208.830 56.100 209.230 ;
        RECT 53.220 206.830 53.540 208.030 ;
        RECT 54.500 207.230 56.740 207.630 ;
        RECT 57.060 206.830 57.380 208.030 ;
        RECT 53.860 205.630 56.100 206.030 ;
        RECT 53.860 201.330 56.100 201.730 ;
        RECT 53.220 199.330 53.540 200.530 ;
        RECT 54.500 199.730 56.740 200.130 ;
        RECT 57.060 199.330 57.380 200.530 ;
        RECT 53.860 198.130 56.100 198.530 ;
        RECT 53.860 194.330 56.100 194.730 ;
        RECT 53.220 192.330 53.540 193.530 ;
        RECT 54.500 192.730 56.740 193.130 ;
        RECT 57.060 192.330 57.380 193.530 ;
        RECT 53.860 191.130 56.100 191.530 ;
        RECT 57.700 190.770 61.900 209.810 ;
        RECT 62.860 208.330 65.100 208.730 ;
        RECT 62.220 206.330 62.540 207.530 ;
        RECT 63.500 206.730 65.740 207.130 ;
        RECT 66.060 206.330 66.380 207.530 ;
        RECT 62.860 205.130 65.100 205.530 ;
        RECT 62.860 201.330 65.100 201.730 ;
        RECT 62.220 199.330 62.540 200.530 ;
        RECT 63.500 199.730 65.740 200.130 ;
        RECT 66.060 199.330 66.380 200.530 ;
        RECT 62.860 198.130 65.100 198.530 ;
        RECT 62.860 194.330 65.100 194.730 ;
        RECT 62.220 192.330 62.540 193.530 ;
        RECT 63.500 192.730 65.740 193.130 ;
        RECT 66.060 192.330 66.380 193.530 ;
        RECT 62.860 191.130 65.100 191.530 ;
        RECT 66.700 190.770 70.900 209.810 ;
        RECT 71.860 208.330 74.100 208.730 ;
        RECT 71.220 206.330 71.540 207.530 ;
        RECT 72.500 206.730 74.740 207.130 ;
        RECT 75.060 206.330 75.380 207.530 ;
        RECT 71.860 205.130 74.100 205.530 ;
        RECT 71.860 201.330 74.100 201.730 ;
        RECT 71.220 199.330 71.540 200.530 ;
        RECT 72.500 199.730 74.740 200.130 ;
        RECT 75.060 199.330 75.380 200.530 ;
        RECT 71.860 198.130 74.100 198.530 ;
        RECT 71.860 194.330 74.100 194.730 ;
        RECT 71.220 192.330 71.540 193.530 ;
        RECT 72.500 192.730 74.740 193.130 ;
        RECT 75.060 192.330 75.380 193.530 ;
        RECT 71.860 191.130 74.100 191.530 ;
        RECT 75.700 190.770 79.900 209.810 ;
        RECT 80.860 208.330 83.100 208.730 ;
        RECT 80.220 206.330 80.540 207.530 ;
        RECT 81.500 206.730 83.740 207.130 ;
        RECT 84.060 206.330 84.380 207.530 ;
        RECT 80.860 205.130 83.100 205.530 ;
        RECT 84.700 202.310 97.900 209.810 ;
        RECT 98.860 208.330 101.100 208.730 ;
        RECT 98.220 206.330 98.540 207.530 ;
        RECT 99.500 206.730 101.740 207.130 ;
        RECT 102.060 206.330 102.380 207.530 ;
        RECT 98.860 205.130 101.100 205.530 ;
        RECT 80.860 201.330 83.100 201.730 ;
        RECT 80.220 199.330 80.540 200.530 ;
        RECT 81.500 199.730 83.740 200.130 ;
        RECT 84.060 199.330 84.380 200.530 ;
        RECT 80.860 198.130 83.100 198.530 ;
        RECT 84.700 197.770 88.900 202.310 ;
        RECT 89.860 201.330 92.100 201.730 ;
        RECT 89.220 199.330 89.540 200.530 ;
        RECT 90.500 199.730 92.740 200.130 ;
        RECT 93.060 199.330 93.380 200.530 ;
        RECT 89.860 198.130 92.100 198.530 ;
        RECT 93.700 197.770 97.900 202.310 ;
        RECT 102.700 202.310 116.300 209.810 ;
        RECT 117.900 208.330 120.140 208.730 ;
        RECT 116.620 206.330 116.940 207.530 ;
        RECT 117.260 206.730 119.500 207.130 ;
        RECT 120.460 206.330 120.780 207.530 ;
        RECT 117.900 205.130 120.140 205.530 ;
        RECT 98.860 201.330 101.100 201.730 ;
        RECT 98.220 199.330 98.540 200.530 ;
        RECT 99.500 199.730 101.740 200.130 ;
        RECT 102.060 199.330 102.380 200.530 ;
        RECT 98.860 198.130 101.100 198.530 ;
        RECT 80.860 194.330 83.100 194.730 ;
        RECT 80.220 192.330 80.540 193.530 ;
        RECT 81.500 192.730 83.740 193.130 ;
        RECT 84.060 192.330 84.380 193.530 ;
        RECT 80.860 191.130 83.100 191.530 ;
        RECT 84.700 190.770 97.900 197.770 ;
        RECT 102.700 197.770 107.300 202.310 ;
        RECT 108.900 201.330 111.140 201.730 ;
        RECT 107.620 199.330 107.940 200.530 ;
        RECT 108.260 199.730 110.500 200.130 ;
        RECT 111.460 199.330 111.780 200.530 ;
        RECT 108.900 198.130 111.140 198.530 ;
        RECT 112.100 197.770 116.300 202.310 ;
        RECT 117.900 201.330 120.140 201.730 ;
        RECT 116.620 199.330 116.940 200.530 ;
        RECT 117.260 199.730 119.500 200.130 ;
        RECT 120.460 199.330 120.780 200.530 ;
        RECT 117.900 198.130 120.140 198.530 ;
        RECT 98.860 194.330 101.100 194.730 ;
        RECT 98.220 192.330 98.540 193.530 ;
        RECT 99.500 192.730 101.740 193.130 ;
        RECT 102.060 192.330 102.380 193.530 ;
        RECT 98.860 191.130 101.100 191.530 ;
        RECT 102.700 190.770 116.300 197.770 ;
        RECT 117.900 194.330 120.140 194.730 ;
        RECT 116.620 192.330 116.940 193.530 ;
        RECT 117.260 192.730 119.500 193.130 ;
        RECT 120.460 192.330 120.780 193.530 ;
        RECT 117.900 191.130 120.140 191.530 ;
        RECT 121.100 190.770 125.300 209.810 ;
        RECT 126.900 208.330 129.140 208.730 ;
        RECT 125.620 206.330 125.940 207.530 ;
        RECT 126.260 206.730 128.500 207.130 ;
        RECT 129.460 206.330 129.780 207.530 ;
        RECT 126.900 205.130 129.140 205.530 ;
        RECT 126.900 201.330 129.140 201.730 ;
        RECT 125.620 199.330 125.940 200.530 ;
        RECT 126.260 199.730 128.500 200.130 ;
        RECT 129.460 199.330 129.780 200.530 ;
        RECT 126.900 198.130 129.140 198.530 ;
        RECT 126.900 194.330 129.140 194.730 ;
        RECT 125.620 192.330 125.940 193.530 ;
        RECT 126.260 192.730 128.500 193.130 ;
        RECT 129.460 192.330 129.780 193.530 ;
        RECT 126.900 191.130 129.140 191.530 ;
        RECT 130.100 190.770 134.300 209.810 ;
        RECT 135.900 208.330 138.140 208.730 ;
        RECT 134.620 206.330 134.940 207.530 ;
        RECT 135.260 206.730 137.500 207.130 ;
        RECT 138.460 206.330 138.780 207.530 ;
        RECT 135.900 205.130 138.140 205.530 ;
        RECT 135.900 201.330 138.140 201.730 ;
        RECT 134.620 199.330 134.940 200.530 ;
        RECT 135.260 199.730 137.500 200.130 ;
        RECT 138.460 199.330 138.780 200.530 ;
        RECT 135.900 198.130 138.140 198.530 ;
        RECT 135.900 194.330 138.140 194.730 ;
        RECT 134.620 192.330 134.940 193.530 ;
        RECT 135.260 192.730 137.500 193.130 ;
        RECT 138.460 192.330 138.780 193.530 ;
        RECT 135.900 191.130 138.140 191.530 ;
        RECT 139.100 190.770 143.300 209.810 ;
        RECT 144.900 208.830 147.140 209.230 ;
        RECT 143.620 206.830 143.940 208.030 ;
        RECT 144.260 207.230 146.500 207.630 ;
        RECT 147.460 206.830 147.780 208.030 ;
        RECT 144.900 205.630 147.140 206.030 ;
        RECT 144.900 201.330 147.140 201.730 ;
        RECT 143.620 199.330 143.940 200.530 ;
        RECT 144.260 199.730 146.500 200.130 ;
        RECT 147.460 199.330 147.780 200.530 ;
        RECT 144.900 198.130 147.140 198.530 ;
        RECT 144.900 194.330 147.140 194.730 ;
        RECT 143.620 192.330 143.940 193.530 ;
        RECT 144.260 192.730 146.500 193.130 ;
        RECT 147.460 192.330 147.780 193.530 ;
        RECT 144.900 191.130 147.140 191.530 ;
        RECT 148.100 190.770 149.060 209.810 ;
        RECT 51.940 189.810 149.060 190.770 ;
        RECT 150.500 194.930 151.140 210.850 ;
        RECT 152.320 208.890 153.760 210.090 ;
        RECT 153.400 205.290 153.760 208.890 ;
        RECT 154.480 208.890 155.920 210.090 ;
        RECT 154.480 205.290 154.840 208.890 ;
        RECT 155.560 205.290 155.920 208.890 ;
        RECT 156.640 208.890 158.080 210.090 ;
        RECT 156.640 205.290 157.000 208.890 ;
        RECT 153.400 195.690 154.840 198.090 ;
        RECT 155.560 195.690 157.000 198.090 ;
        RECT 159.260 194.930 160.500 210.850 ;
        RECT 150.500 192.850 160.500 194.930 ;
        RECT 85.000 189.790 97.500 189.810 ;
        RECT 103.000 189.790 115.500 189.810 ;
        RECT 54.500 187.790 77.000 188.790 ;
        RECT 54.500 171.930 55.140 187.790 ;
        RECT 56.320 185.890 57.760 187.090 ;
        RECT 57.400 182.290 57.760 185.890 ;
        RECT 58.480 185.890 59.920 187.090 ;
        RECT 58.480 182.290 58.840 185.890 ;
        RECT 59.560 182.290 59.920 185.890 ;
        RECT 60.640 185.890 62.080 187.090 ;
        RECT 60.640 182.290 61.000 185.890 ;
        RECT 61.720 182.290 62.080 185.890 ;
        RECT 62.800 185.890 64.240 187.090 ;
        RECT 62.800 182.290 63.160 185.890 ;
        RECT 63.880 182.290 64.240 185.890 ;
        RECT 64.960 185.890 66.400 187.090 ;
        RECT 64.960 182.290 65.320 185.890 ;
        RECT 66.040 182.290 66.400 185.890 ;
        RECT 67.120 185.890 68.560 187.090 ;
        RECT 67.120 182.290 67.480 185.890 ;
        RECT 68.200 182.290 68.560 185.890 ;
        RECT 69.280 185.890 70.720 187.090 ;
        RECT 69.280 182.290 69.640 185.890 ;
        RECT 70.360 182.290 70.720 185.890 ;
        RECT 71.440 185.890 72.880 187.090 ;
        RECT 71.440 182.290 71.800 185.890 ;
        RECT 72.520 182.290 72.880 185.890 ;
        RECT 73.600 185.890 75.040 187.090 ;
        RECT 73.600 182.290 73.960 185.890 ;
        RECT 57.400 172.690 58.840 175.090 ;
        RECT 59.560 172.690 61.000 175.090 ;
        RECT 61.720 172.690 63.160 175.090 ;
        RECT 63.880 172.690 65.320 175.090 ;
        RECT 66.040 172.690 67.480 175.090 ;
        RECT 68.200 172.690 69.640 175.090 ;
        RECT 70.360 172.690 71.800 175.090 ;
        RECT 72.520 172.690 73.960 175.090 ;
        RECT 76.220 172.770 77.000 187.790 ;
        RECT 124.220 188.290 146.420 188.410 ;
        RECT 150.500 188.290 151.140 192.850 ;
        RECT 152.320 190.890 153.760 192.090 ;
        RECT 124.220 187.850 151.140 188.290 ;
        RECT 78.940 186.810 94.660 187.770 ;
        RECT 78.940 174.770 79.900 186.810 ;
        RECT 80.860 185.830 83.100 186.230 ;
        RECT 80.220 183.830 80.540 185.030 ;
        RECT 81.500 184.230 83.740 184.630 ;
        RECT 84.060 183.830 84.380 185.030 ;
        RECT 80.860 182.630 83.100 183.030 ;
        RECT 80.860 178.330 83.100 178.730 ;
        RECT 80.220 176.330 80.540 177.530 ;
        RECT 81.500 176.730 83.740 177.130 ;
        RECT 84.060 176.330 84.380 177.530 ;
        RECT 80.860 175.130 83.100 175.530 ;
        RECT 84.700 174.770 88.900 186.810 ;
        RECT 89.860 185.330 92.100 185.730 ;
        RECT 89.220 183.330 89.540 184.530 ;
        RECT 90.500 183.730 92.740 184.130 ;
        RECT 93.060 183.330 93.380 184.530 ;
        RECT 89.860 182.130 92.100 182.530 ;
        RECT 89.860 178.330 92.100 178.730 ;
        RECT 89.220 176.330 89.540 177.530 ;
        RECT 90.500 176.730 92.740 177.130 ;
        RECT 93.060 176.330 93.380 177.530 ;
        RECT 89.860 175.130 92.100 175.530 ;
        RECT 93.700 174.770 94.660 186.810 ;
        RECT 78.940 173.810 94.660 174.770 ;
        RECT 106.340 186.810 122.060 187.770 ;
        RECT 106.340 174.770 107.300 186.810 ;
        RECT 108.900 185.330 111.140 185.730 ;
        RECT 107.620 183.330 107.940 184.530 ;
        RECT 108.260 183.730 110.500 184.130 ;
        RECT 111.460 183.330 111.780 184.530 ;
        RECT 108.900 182.130 111.140 182.530 ;
        RECT 108.900 178.330 111.140 178.730 ;
        RECT 107.620 176.330 107.940 177.530 ;
        RECT 108.260 176.730 110.500 177.130 ;
        RECT 111.460 176.330 111.780 177.530 ;
        RECT 108.900 175.130 111.140 175.530 ;
        RECT 112.100 174.770 116.300 186.810 ;
        RECT 117.900 185.830 120.140 186.230 ;
        RECT 116.620 183.830 116.940 185.030 ;
        RECT 117.260 184.230 119.500 184.630 ;
        RECT 120.460 183.830 120.780 185.030 ;
        RECT 117.900 182.630 120.140 183.030 ;
        RECT 117.900 178.330 120.140 178.730 ;
        RECT 116.620 176.330 116.940 177.530 ;
        RECT 117.260 176.730 119.500 177.130 ;
        RECT 120.460 176.330 120.780 177.530 ;
        RECT 117.900 175.130 120.140 175.530 ;
        RECT 121.100 174.770 122.060 186.810 ;
        RECT 106.340 173.810 122.060 174.770 ;
        RECT 76.220 172.290 122.060 172.770 ;
        RECT 124.220 172.290 124.780 187.850 ;
        RECT 125.960 185.890 127.400 187.090 ;
        RECT 127.040 182.290 127.400 185.890 ;
        RECT 128.120 185.890 129.560 187.090 ;
        RECT 128.120 182.290 128.480 185.890 ;
        RECT 129.200 182.290 129.560 185.890 ;
        RECT 130.280 185.890 131.720 187.090 ;
        RECT 130.280 182.290 130.640 185.890 ;
        RECT 131.360 182.290 131.720 185.890 ;
        RECT 132.440 185.890 133.880 187.090 ;
        RECT 132.440 182.290 132.800 185.890 ;
        RECT 133.520 182.290 133.880 185.890 ;
        RECT 134.600 185.890 136.040 187.090 ;
        RECT 134.600 182.290 134.960 185.890 ;
        RECT 135.680 182.290 136.040 185.890 ;
        RECT 136.760 185.890 138.200 187.090 ;
        RECT 136.760 182.290 137.120 185.890 ;
        RECT 137.840 182.290 138.200 185.890 ;
        RECT 138.920 185.890 140.360 187.090 ;
        RECT 138.920 182.290 139.280 185.890 ;
        RECT 140.000 182.290 140.360 185.890 ;
        RECT 141.080 185.890 142.520 187.090 ;
        RECT 141.080 182.290 141.440 185.890 ;
        RECT 142.160 182.290 142.520 185.890 ;
        RECT 143.240 185.890 144.680 187.090 ;
        RECT 143.240 182.290 143.600 185.890 ;
        RECT 145.860 176.930 151.140 187.850 ;
        RECT 153.400 187.290 153.760 190.890 ;
        RECT 154.480 190.890 155.920 192.090 ;
        RECT 154.480 187.290 154.840 190.890 ;
        RECT 155.560 187.290 155.920 190.890 ;
        RECT 156.640 190.890 158.080 192.090 ;
        RECT 156.640 187.290 157.000 190.890 ;
        RECT 153.400 177.690 154.840 180.090 ;
        RECT 155.560 177.690 157.000 180.090 ;
        RECT 159.260 176.930 160.500 192.850 ;
        RECT 127.040 172.690 128.480 175.090 ;
        RECT 129.200 172.690 130.640 175.090 ;
        RECT 131.360 172.690 132.800 175.090 ;
        RECT 133.520 172.690 134.960 175.090 ;
        RECT 135.680 172.690 137.120 175.090 ;
        RECT 137.840 172.690 139.280 175.090 ;
        RECT 140.000 172.690 141.440 175.090 ;
        RECT 142.160 172.690 143.600 175.090 ;
        RECT 145.860 174.850 160.500 176.930 ;
        RECT 76.220 171.930 124.780 172.290 ;
        RECT 145.860 171.930 151.140 174.850 ;
        RECT 152.320 172.890 153.760 174.090 ;
        RECT 54.500 171.810 151.140 171.930 ;
        RECT 54.500 169.850 79.900 171.810 ;
        RECT 80.860 170.330 83.100 170.730 ;
        RECT 16.990 151.180 17.890 167.230 ;
        RECT 22.690 166.780 22.990 167.680 ;
        RECT 20.590 166.480 24.190 166.780 ;
        RECT 18.790 166.080 19.690 166.380 ;
        RECT 25.090 166.080 25.990 166.380 ;
        RECT 19.390 165.780 20.290 166.080 ;
        RECT 18.790 165.280 19.690 165.580 ;
        RECT 19.990 165.480 20.290 165.780 ;
        RECT 20.590 165.980 21.430 166.000 ;
        RECT 23.290 165.980 24.130 166.000 ;
        RECT 20.590 165.680 21.490 165.980 ;
        RECT 23.290 165.680 24.190 165.980 ;
        RECT 19.000 164.980 19.300 165.280 ;
        RECT 19.990 165.180 20.890 165.480 ;
        RECT 25.090 165.280 25.990 165.580 ;
        RECT 19.000 164.680 19.870 164.980 ;
        RECT 20.590 164.880 24.190 165.180 ;
        RECT 21.820 164.380 22.430 164.400 ;
        RECT 20.590 164.080 24.190 164.380 ;
        RECT 18.790 163.680 19.690 163.980 ;
        RECT 25.090 163.680 25.990 163.980 ;
        RECT 19.390 163.380 20.290 163.680 ;
        RECT 18.790 162.880 19.690 163.180 ;
        RECT 19.990 163.080 20.290 163.380 ;
        RECT 20.590 163.580 21.430 163.600 ;
        RECT 23.290 163.580 24.130 163.600 ;
        RECT 20.590 163.280 21.490 163.580 ;
        RECT 23.290 163.280 24.190 163.580 ;
        RECT 19.990 162.780 20.890 163.080 ;
        RECT 25.090 162.880 25.990 163.180 ;
        RECT 20.590 162.480 24.190 162.780 ;
        RECT 25.550 162.260 25.870 162.880 ;
        RECT 20.060 161.680 21.490 161.980 ;
        RECT 23.290 161.680 24.790 161.980 ;
        RECT 24.490 161.580 24.790 161.680 ;
        RECT 18.790 161.280 19.690 161.580 ;
        RECT 24.490 161.280 25.990 161.580 ;
        RECT 20.590 161.180 21.430 161.200 ;
        RECT 23.290 161.180 24.130 161.200 ;
        RECT 20.590 160.880 21.490 161.180 ;
        RECT 23.290 160.880 24.190 161.180 ;
        RECT 18.820 160.400 20.240 160.700 ;
        RECT 19.940 160.380 20.240 160.400 ;
        RECT 19.940 160.080 24.190 160.380 ;
        RECT 18.790 159.680 19.690 159.980 ;
        RECT 25.090 159.680 25.990 159.980 ;
        RECT 19.390 159.380 20.290 159.680 ;
        RECT 18.790 158.880 19.690 159.180 ;
        RECT 19.990 159.080 20.290 159.380 ;
        RECT 20.590 159.580 21.430 159.600 ;
        RECT 23.290 159.580 24.130 159.600 ;
        RECT 20.590 159.280 21.490 159.580 ;
        RECT 23.290 159.280 24.190 159.580 ;
        RECT 19.040 157.580 19.340 158.880 ;
        RECT 19.990 158.780 20.890 159.080 ;
        RECT 25.090 158.880 25.990 159.180 ;
        RECT 20.590 158.480 24.190 158.780 ;
        RECT 20.590 157.980 21.430 158.000 ;
        RECT 20.590 157.680 21.490 157.980 ;
        RECT 21.790 157.680 24.190 157.980 ;
        RECT 18.790 157.280 19.690 157.580 ;
        RECT 21.790 157.180 22.090 157.680 ;
        RECT 25.325 157.580 25.660 158.305 ;
        RECT 25.090 157.280 25.990 157.580 ;
        RECT 19.970 156.880 22.090 157.180 ;
        RECT 23.290 156.880 24.190 157.180 ;
        RECT 19.360 156.780 19.660 156.800 ;
        RECT 18.790 156.480 19.690 156.780 ;
        RECT 25.090 156.480 25.990 156.780 ;
        RECT 19.360 156.160 19.660 156.480 ;
        RECT 20.590 156.380 21.430 156.400 ;
        RECT 23.290 156.380 24.130 156.400 ;
        RECT 19.360 155.860 20.420 156.160 ;
        RECT 20.590 156.080 21.490 156.380 ;
        RECT 23.290 156.080 24.190 156.380 ;
        RECT 20.120 155.580 20.420 155.860 ;
        RECT 20.120 155.280 24.190 155.580 ;
        RECT 18.790 154.880 19.690 155.180 ;
        RECT 25.090 154.880 25.990 155.180 ;
        RECT 19.150 154.500 19.450 154.880 ;
        RECT 20.590 154.780 21.430 154.800 ;
        RECT 23.290 154.780 24.130 154.800 ;
        RECT 19.150 154.200 20.310 154.500 ;
        RECT 20.590 154.480 21.490 154.780 ;
        RECT 23.290 154.480 24.190 154.780 ;
        RECT 20.010 153.980 20.310 154.200 ;
        RECT 24.400 154.090 25.870 154.390 ;
        RECT 24.400 153.980 24.700 154.090 ;
        RECT 20.010 153.680 24.700 153.980 ;
        RECT 18.790 153.280 19.690 153.580 ;
        RECT 25.090 153.280 25.990 153.580 ;
        RECT 19.390 152.980 20.290 153.280 ;
        RECT 18.790 152.480 19.690 152.780 ;
        RECT 19.990 152.680 20.290 152.980 ;
        RECT 20.590 153.180 21.430 153.200 ;
        RECT 23.290 153.180 24.130 153.200 ;
        RECT 20.590 152.880 21.490 153.180 ;
        RECT 23.290 152.880 24.190 153.180 ;
        RECT 19.990 152.380 20.890 152.680 ;
        RECT 25.090 152.480 25.990 152.780 ;
        RECT 20.590 152.080 24.190 152.380 ;
        RECT 20.590 151.580 21.430 151.600 ;
        RECT 23.290 151.580 24.130 151.600 ;
        RECT 19.990 151.280 21.490 151.580 ;
        RECT 23.290 151.280 24.790 151.580 ;
        RECT 19.990 151.180 20.290 151.280 ;
        RECT 16.990 150.880 20.290 151.180 ;
        RECT 16.990 150.030 17.890 150.880 ;
        RECT 19.990 150.780 20.290 150.880 ;
        RECT 24.490 151.180 24.790 151.280 ;
        RECT 26.890 151.180 27.790 167.230 ;
        RECT 24.490 150.880 27.790 151.180 ;
        RECT 20.590 150.780 21.430 150.800 ;
        RECT 23.290 150.780 24.130 150.800 ;
        RECT 24.490 150.780 24.790 150.880 ;
        RECT 19.990 150.480 21.490 150.780 ;
        RECT 23.290 150.480 24.790 150.780 ;
        RECT 26.890 150.030 27.790 150.880 ;
        RECT 54.500 153.930 55.140 169.850 ;
        RECT 73.840 169.090 75.040 169.850 ;
        RECT 56.320 167.890 57.760 169.090 ;
        RECT 57.400 164.290 57.760 167.890 ;
        RECT 58.480 167.890 59.920 169.090 ;
        RECT 58.480 164.290 58.840 167.890 ;
        RECT 59.560 164.290 59.920 167.890 ;
        RECT 60.640 167.890 62.080 169.090 ;
        RECT 60.640 164.290 61.000 167.890 ;
        RECT 61.720 164.290 62.080 167.890 ;
        RECT 62.800 167.890 64.240 169.090 ;
        RECT 62.800 164.290 63.160 167.890 ;
        RECT 63.880 164.290 64.240 167.890 ;
        RECT 64.960 167.890 66.400 169.090 ;
        RECT 64.960 164.290 65.320 167.890 ;
        RECT 66.040 164.290 66.400 167.890 ;
        RECT 67.120 167.890 68.560 169.090 ;
        RECT 67.120 164.290 67.480 167.890 ;
        RECT 68.200 164.290 68.560 167.890 ;
        RECT 69.280 167.890 70.720 169.090 ;
        RECT 69.280 164.290 69.640 167.890 ;
        RECT 70.360 164.290 70.720 167.890 ;
        RECT 71.440 167.890 72.880 169.090 ;
        RECT 71.440 164.290 71.800 167.890 ;
        RECT 72.520 164.290 72.880 167.890 ;
        RECT 73.600 167.890 75.040 169.090 ;
        RECT 73.600 164.290 73.960 167.890 ;
        RECT 76.220 161.790 79.900 169.850 ;
        RECT 80.220 168.330 80.540 169.530 ;
        RECT 81.500 168.730 83.740 169.130 ;
        RECT 84.060 168.330 84.380 169.530 ;
        RECT 80.860 167.130 83.100 167.530 ;
        RECT 80.860 165.330 83.100 165.730 ;
        RECT 80.220 163.330 80.540 164.530 ;
        RECT 81.500 163.730 83.740 164.130 ;
        RECT 84.060 163.330 84.380 164.530 ;
        RECT 80.860 162.130 83.100 162.530 ;
        RECT 84.700 161.790 88.900 171.810 ;
        RECT 89.860 170.330 92.100 170.730 ;
        RECT 89.220 168.330 89.540 169.530 ;
        RECT 90.500 168.730 92.740 169.130 ;
        RECT 93.060 168.330 93.380 169.530 ;
        RECT 89.860 167.130 92.100 167.530 ;
        RECT 89.860 165.330 92.100 165.730 ;
        RECT 89.220 163.330 89.540 164.530 ;
        RECT 90.500 163.730 92.740 164.130 ;
        RECT 93.060 163.330 93.380 164.530 ;
        RECT 89.860 162.130 92.100 162.530 ;
        RECT 93.700 161.790 107.300 171.810 ;
        RECT 108.900 170.330 111.140 170.730 ;
        RECT 107.620 168.330 107.940 169.530 ;
        RECT 108.260 168.730 110.500 169.130 ;
        RECT 111.460 168.330 111.780 169.530 ;
        RECT 108.900 167.130 111.140 167.530 ;
        RECT 108.900 165.330 111.140 165.730 ;
        RECT 107.620 163.330 107.940 164.530 ;
        RECT 108.260 163.730 110.500 164.130 ;
        RECT 111.460 163.330 111.780 164.530 ;
        RECT 108.900 162.130 111.140 162.530 ;
        RECT 76.220 161.770 107.300 161.790 ;
        RECT 112.100 161.770 116.300 171.810 ;
        RECT 117.900 170.330 120.140 170.730 ;
        RECT 121.100 169.850 151.140 171.810 ;
        RECT 116.620 168.330 116.940 169.530 ;
        RECT 117.260 168.730 119.500 169.130 ;
        RECT 120.460 168.330 120.780 169.530 ;
        RECT 117.900 167.130 120.140 167.530 ;
        RECT 117.900 165.330 120.140 165.730 ;
        RECT 116.620 163.330 116.940 164.530 ;
        RECT 117.260 163.730 119.500 164.130 ;
        RECT 120.460 163.330 120.780 164.530 ;
        RECT 117.900 162.130 120.140 162.530 ;
        RECT 121.100 161.770 124.780 169.850 ;
        RECT 125.960 169.090 127.160 169.850 ;
        RECT 125.960 167.890 127.400 169.090 ;
        RECT 127.040 164.290 127.400 167.890 ;
        RECT 128.120 167.890 129.560 169.090 ;
        RECT 128.120 164.290 128.480 167.890 ;
        RECT 129.200 164.290 129.560 167.890 ;
        RECT 130.280 167.890 131.720 169.090 ;
        RECT 130.280 164.290 130.640 167.890 ;
        RECT 131.360 164.290 131.720 167.890 ;
        RECT 132.440 167.890 133.880 169.090 ;
        RECT 132.440 164.290 132.800 167.890 ;
        RECT 133.520 164.290 133.880 167.890 ;
        RECT 134.600 167.890 136.040 169.090 ;
        RECT 134.600 164.290 134.960 167.890 ;
        RECT 135.680 164.290 136.040 167.890 ;
        RECT 136.760 167.890 138.200 169.090 ;
        RECT 136.760 164.290 137.120 167.890 ;
        RECT 137.840 164.290 138.200 167.890 ;
        RECT 138.920 167.890 140.360 169.090 ;
        RECT 138.920 164.290 139.280 167.890 ;
        RECT 140.000 164.290 140.360 167.890 ;
        RECT 141.080 167.890 142.520 169.090 ;
        RECT 141.080 164.290 141.440 167.890 ;
        RECT 142.160 164.290 142.520 167.890 ;
        RECT 143.240 167.890 144.680 169.090 ;
        RECT 143.240 164.290 143.600 167.890 ;
        RECT 76.220 160.810 124.780 161.770 ;
        RECT 76.220 160.290 107.000 160.810 ;
        RECT 57.400 154.690 58.840 157.090 ;
        RECT 59.560 154.690 61.000 157.090 ;
        RECT 61.720 154.690 63.160 157.090 ;
        RECT 63.880 154.690 65.320 157.090 ;
        RECT 66.040 154.690 67.480 157.090 ;
        RECT 68.200 154.690 69.640 157.090 ;
        RECT 70.360 154.690 71.800 157.090 ;
        RECT 72.520 154.690 73.960 157.090 ;
        RECT 76.220 156.685 102.500 160.290 ;
        RECT 104.600 157.670 105.500 158.890 ;
        RECT 107.450 158.140 111.800 158.440 ;
        RECT 106.400 157.740 107.300 158.040 ;
        RECT 112.700 157.740 113.600 158.040 ;
        RECT 103.420 156.710 105.500 157.670 ;
        RECT 108.260 157.640 109.100 157.660 ;
        RECT 110.960 157.640 111.800 157.660 ;
        RECT 108.200 157.340 109.100 157.640 ;
        RECT 110.900 157.340 111.800 157.640 ;
        RECT 112.100 157.440 113.000 157.740 ;
        RECT 114.500 157.630 115.400 158.890 ;
        RECT 106.400 156.940 107.300 157.240 ;
        RECT 112.100 157.140 112.400 157.440 ;
        RECT 111.500 156.840 112.400 157.140 ;
        RECT 112.700 156.940 114.050 157.240 ;
        RECT 76.220 153.930 80.805 156.685 ;
        RECT 54.500 152.595 80.805 153.930 ;
        RECT 81.115 152.905 84.585 156.375 ;
        RECT 84.895 152.595 88.805 156.685 ;
        RECT 89.115 152.905 92.585 156.375 ;
        RECT 92.895 152.595 96.805 156.685 ;
        RECT 97.115 152.905 100.585 156.375 ;
        RECT 100.895 154.290 102.500 156.685 ;
        RECT 104.600 156.090 105.500 156.710 ;
        RECT 108.200 156.540 111.800 156.840 ;
        RECT 114.500 156.750 116.640 157.630 ;
        RECT 114.500 156.090 115.400 156.750 ;
        RECT 115.760 155.350 116.640 156.750 ;
        RECT 100.895 153.790 104.500 154.290 ;
        RECT 100.895 152.595 104.700 153.790 ;
        RECT 109.350 153.340 109.650 153.940 ;
        RECT 122.000 153.930 124.780 160.810 ;
        RECT 145.860 158.930 151.140 169.850 ;
        RECT 153.400 169.290 153.760 172.890 ;
        RECT 154.480 172.890 155.920 174.090 ;
        RECT 154.480 169.290 154.840 172.890 ;
        RECT 155.560 169.290 155.920 172.890 ;
        RECT 156.640 172.890 158.080 174.090 ;
        RECT 156.640 169.290 157.000 172.890 ;
        RECT 153.400 159.690 154.840 162.090 ;
        RECT 155.560 159.690 157.000 162.090 ;
        RECT 159.260 158.930 160.500 174.850 ;
        RECT 127.040 154.690 128.480 157.090 ;
        RECT 129.200 154.690 130.640 157.090 ;
        RECT 131.360 154.690 132.800 157.090 ;
        RECT 133.520 154.690 134.960 157.090 ;
        RECT 135.680 154.690 137.120 157.090 ;
        RECT 137.840 154.690 139.280 157.090 ;
        RECT 140.000 154.690 141.440 157.090 ;
        RECT 142.160 154.690 143.600 157.090 ;
        RECT 145.860 156.850 160.500 158.930 ;
        RECT 145.860 156.090 151.140 156.850 ;
        RECT 145.860 154.890 153.760 156.090 ;
        RECT 145.860 153.930 151.140 154.890 ;
        RECT 110.100 153.340 110.940 153.360 ;
        RECT 107.400 153.040 111.000 153.340 ;
        RECT 105.600 152.640 107.100 152.940 ;
        RECT 111.900 152.640 112.800 152.940 ;
        RECT 54.500 151.790 104.700 152.595 ;
        RECT 9.720 139.940 13.700 139.950 ;
        RECT 9.720 138.010 44.165 139.940 ;
        RECT 42.235 135.915 44.165 138.010 ;
        RECT 54.500 135.930 55.140 151.790 ;
        RECT 56.320 149.890 57.760 151.090 ;
        RECT 57.400 146.290 57.760 149.890 ;
        RECT 58.480 149.890 59.920 151.090 ;
        RECT 58.480 146.290 58.840 149.890 ;
        RECT 59.560 146.290 59.920 149.890 ;
        RECT 60.640 149.890 62.080 151.090 ;
        RECT 60.640 146.290 61.000 149.890 ;
        RECT 61.720 146.290 62.080 149.890 ;
        RECT 62.800 149.890 64.240 151.090 ;
        RECT 62.800 146.290 63.160 149.890 ;
        RECT 63.880 146.290 64.240 149.890 ;
        RECT 64.960 149.890 66.400 151.090 ;
        RECT 64.960 146.290 65.320 149.890 ;
        RECT 66.040 146.290 66.400 149.890 ;
        RECT 67.120 149.890 68.560 151.090 ;
        RECT 67.120 146.290 67.480 149.890 ;
        RECT 68.200 146.290 68.560 149.890 ;
        RECT 69.280 149.890 70.720 151.090 ;
        RECT 69.280 146.290 69.640 149.890 ;
        RECT 70.360 146.290 70.720 149.890 ;
        RECT 71.440 149.890 72.880 151.090 ;
        RECT 71.440 146.290 71.800 149.890 ;
        RECT 72.520 146.290 72.880 149.890 ;
        RECT 73.600 149.890 75.040 151.090 ;
        RECT 73.600 146.290 73.960 149.890 ;
        RECT 76.220 148.685 104.700 151.790 ;
        RECT 106.800 151.740 107.100 152.640 ;
        RECT 107.400 152.540 108.240 152.560 ;
        RECT 110.100 152.540 110.940 152.560 ;
        RECT 107.400 152.240 108.300 152.540 ;
        RECT 110.100 152.240 111.000 152.540 ;
        RECT 107.400 151.740 108.240 151.760 ;
        RECT 106.800 151.440 111.000 151.740 ;
        RECT 105.600 151.340 106.440 151.360 ;
        RECT 105.600 151.040 106.500 151.340 ;
        RECT 111.300 151.040 112.800 151.340 ;
        RECT 107.400 150.640 111.000 150.940 ;
        RECT 105.600 150.240 106.500 150.540 ;
        RECT 107.400 149.840 108.300 150.140 ;
        RECT 105.600 149.740 106.440 149.760 ;
        RECT 105.600 149.440 106.500 149.740 ;
        RECT 107.400 149.340 108.240 149.360 ;
        RECT 109.500 149.340 109.800 150.640 ;
        RECT 110.100 150.140 110.940 150.160 ;
        RECT 110.100 149.840 111.000 150.140 ;
        RECT 107.400 149.040 108.300 149.340 ;
        RECT 109.500 149.040 111.000 149.340 ;
        RECT 76.220 144.595 80.805 148.685 ;
        RECT 81.115 144.905 84.585 148.375 ;
        RECT 84.895 144.595 88.805 148.685 ;
        RECT 89.115 144.905 92.585 148.375 ;
        RECT 92.895 144.595 96.805 148.685 ;
        RECT 97.115 144.905 100.585 148.375 ;
        RECT 100.895 144.595 104.700 148.685 ;
        RECT 107.400 148.540 108.240 148.560 ;
        RECT 107.400 148.240 111.000 148.540 ;
        RECT 105.600 147.840 106.500 148.140 ;
        RECT 106.200 147.540 107.100 147.840 ;
        RECT 105.600 147.040 106.500 147.340 ;
        RECT 105.600 145.740 106.440 145.760 ;
        RECT 105.600 145.440 106.500 145.740 ;
        RECT 76.220 140.685 104.700 144.595 ;
        RECT 106.800 144.140 107.100 147.540 ;
        RECT 107.400 147.440 108.300 147.740 ;
        RECT 110.100 147.440 111.000 147.740 ;
        RECT 107.400 146.940 108.240 146.960 ;
        RECT 110.100 146.940 110.940 146.960 ;
        RECT 107.400 146.640 108.300 146.940 ;
        RECT 110.100 146.640 111.000 146.940 ;
        RECT 110.100 146.140 110.940 146.160 ;
        RECT 107.400 145.840 111.000 146.140 ;
        RECT 107.400 145.340 108.240 145.360 ;
        RECT 110.100 145.340 110.940 145.360 ;
        RECT 107.400 145.040 108.300 145.340 ;
        RECT 110.100 145.040 111.000 145.340 ;
        RECT 107.400 144.540 108.240 144.560 ;
        RECT 107.400 144.240 111.000 144.540 ;
        RECT 105.600 143.840 107.100 144.140 ;
        RECT 105.600 143.040 106.500 143.340 ;
        RECT 105.600 141.740 106.440 141.760 ;
        RECT 105.600 141.440 106.500 141.740 ;
        RECT 57.400 136.690 58.840 139.090 ;
        RECT 59.560 136.690 61.000 139.090 ;
        RECT 61.720 136.690 63.160 139.090 ;
        RECT 63.880 136.690 65.320 139.090 ;
        RECT 66.040 136.690 67.480 139.090 ;
        RECT 68.200 136.690 69.640 139.090 ;
        RECT 70.360 136.690 71.800 139.090 ;
        RECT 72.520 136.690 73.960 139.090 ;
        RECT 76.220 136.595 80.805 140.685 ;
        RECT 81.115 136.905 84.585 140.375 ;
        RECT 84.895 136.595 88.805 140.685 ;
        RECT 89.115 136.905 92.585 140.375 ;
        RECT 92.895 136.595 96.805 140.685 ;
        RECT 97.115 136.905 100.585 140.375 ;
        RECT 100.895 136.595 104.700 140.685 ;
        RECT 105.600 140.640 106.500 140.940 ;
        RECT 106.800 139.740 107.100 143.840 ;
        RECT 107.400 143.440 108.300 143.740 ;
        RECT 107.400 142.940 108.240 142.960 ;
        RECT 107.400 142.640 108.300 142.940 ;
        RECT 108.600 142.140 108.900 144.240 ;
        RECT 110.100 143.440 111.000 143.740 ;
        RECT 110.100 142.940 110.940 142.960 ;
        RECT 110.100 142.640 111.000 142.940 ;
        RECT 107.400 141.840 111.000 142.140 ;
        RECT 111.300 141.740 111.600 151.040 ;
        RECT 111.900 150.540 112.740 150.560 ;
        RECT 111.900 150.240 112.800 150.540 ;
        RECT 111.900 149.440 112.800 149.740 ;
        RECT 111.900 148.140 112.740 148.160 ;
        RECT 111.900 147.840 112.800 148.140 ;
        RECT 111.900 147.340 112.740 147.360 ;
        RECT 111.900 147.040 112.800 147.340 ;
        RECT 111.900 145.440 112.800 145.740 ;
        RECT 111.900 144.140 112.740 144.160 ;
        RECT 111.900 143.840 112.800 144.140 ;
        RECT 111.900 143.340 112.740 143.360 ;
        RECT 111.900 143.040 112.800 143.340 ;
        RECT 111.300 141.440 112.800 141.740 ;
        RECT 107.400 141.040 108.300 141.340 ;
        RECT 110.100 141.040 111.000 141.340 ;
        RECT 107.400 140.540 108.240 140.560 ;
        RECT 110.100 140.540 110.940 140.560 ;
        RECT 107.400 140.240 108.300 140.540 ;
        RECT 110.100 140.240 111.000 140.540 ;
        RECT 111.300 139.740 111.600 141.440 ;
        RECT 111.900 140.640 112.800 140.940 ;
        RECT 112.350 140.140 112.650 140.640 ;
        RECT 106.800 139.440 111.600 139.740 ;
        RECT 105.600 139.040 106.500 139.340 ;
        RECT 111.900 139.040 112.800 139.340 ;
        RECT 107.400 138.940 108.240 138.960 ;
        RECT 110.100 138.940 110.940 138.960 ;
        RECT 107.400 138.640 108.300 138.940 ;
        RECT 110.100 138.640 111.000 138.940 ;
        RECT 111.300 138.740 112.200 139.040 ;
        RECT 107.400 138.140 108.240 138.160 ;
        RECT 110.100 138.140 110.940 138.160 ;
        RECT 107.400 137.840 108.900 138.140 ;
        RECT 110.100 137.840 111.000 138.140 ;
        RECT 105.600 137.740 106.440 137.760 ;
        RECT 105.600 137.440 106.500 137.740 ;
        RECT 108.600 137.340 108.900 137.840 ;
        RECT 110.100 137.340 110.940 137.360 ;
        RECT 111.300 137.340 111.600 138.740 ;
        RECT 111.900 137.440 112.800 137.740 ;
        RECT 107.400 137.040 108.300 137.340 ;
        RECT 108.600 137.040 111.600 137.340 ;
        RECT 105.350 136.640 106.500 136.940 ;
        RECT 111.900 136.640 112.800 136.940 ;
        RECT 76.220 135.930 104.700 136.595 ;
        RECT 105.790 135.940 106.090 136.640 ;
        RECT 107.400 136.540 108.240 136.560 ;
        RECT 110.100 136.540 110.940 136.560 ;
        RECT 107.400 136.240 108.300 136.540 ;
        RECT 110.100 136.240 111.000 136.540 ;
        RECT 54.500 135.915 104.700 135.930 ;
        RECT 42.235 135.340 104.700 135.915 ;
        RECT 107.400 135.740 108.240 135.760 ;
        RECT 110.100 135.740 110.940 135.760 ;
        RECT 106.800 135.440 108.300 135.740 ;
        RECT 110.100 135.440 111.600 135.740 ;
        RECT 106.800 135.340 107.100 135.440 ;
        RECT 42.235 135.040 107.100 135.340 ;
        RECT 42.235 134.190 104.700 135.040 ;
        RECT 106.800 134.940 107.100 135.040 ;
        RECT 111.300 135.340 111.600 135.440 ;
        RECT 113.700 135.340 114.600 153.790 ;
        RECT 122.000 153.290 151.140 153.930 ;
        RECT 111.300 135.040 114.600 135.340 ;
        RECT 107.400 134.940 108.240 134.960 ;
        RECT 110.100 134.940 110.940 134.960 ;
        RECT 111.300 134.940 111.600 135.040 ;
        RECT 106.800 134.640 108.300 134.940 ;
        RECT 110.100 134.640 111.600 134.940 ;
        RECT 42.235 133.985 104.500 134.190 ;
        RECT 54.500 133.790 104.500 133.985 ;
        RECT 54.500 117.930 55.140 133.790 ;
        RECT 56.320 131.890 57.760 133.090 ;
        RECT 57.400 128.290 57.760 131.890 ;
        RECT 58.480 131.890 59.920 133.090 ;
        RECT 58.480 128.290 58.840 131.890 ;
        RECT 59.560 128.290 59.920 131.890 ;
        RECT 60.640 131.890 62.080 133.090 ;
        RECT 60.640 128.290 61.000 131.890 ;
        RECT 61.720 128.290 62.080 131.890 ;
        RECT 62.800 131.890 64.240 133.090 ;
        RECT 62.800 128.290 63.160 131.890 ;
        RECT 63.880 128.290 64.240 131.890 ;
        RECT 64.960 131.890 66.400 133.090 ;
        RECT 64.960 128.290 65.320 131.890 ;
        RECT 66.040 128.290 66.400 131.890 ;
        RECT 67.120 131.890 68.560 133.090 ;
        RECT 67.120 128.290 67.480 131.890 ;
        RECT 68.200 128.290 68.560 131.890 ;
        RECT 69.280 131.890 70.720 133.090 ;
        RECT 69.280 128.290 69.640 131.890 ;
        RECT 70.360 128.290 70.720 131.890 ;
        RECT 71.440 131.890 72.880 133.090 ;
        RECT 71.440 128.290 71.800 131.890 ;
        RECT 72.520 128.290 72.880 131.890 ;
        RECT 73.600 131.890 75.040 133.090 ;
        RECT 73.600 128.290 73.960 131.890 ;
        RECT 57.400 118.690 58.840 121.090 ;
        RECT 59.560 118.690 61.000 121.090 ;
        RECT 61.720 118.690 63.160 121.090 ;
        RECT 63.880 118.690 65.320 121.090 ;
        RECT 66.040 118.690 67.480 121.090 ;
        RECT 68.200 118.690 69.640 121.090 ;
        RECT 70.360 118.690 71.800 121.090 ;
        RECT 72.520 118.690 73.960 121.090 ;
        RECT 76.220 117.930 79.140 133.790 ;
        RECT 80.320 131.890 81.760 133.090 ;
        RECT 81.400 128.290 81.760 131.890 ;
        RECT 82.480 131.890 83.920 133.090 ;
        RECT 82.480 128.290 82.840 131.890 ;
        RECT 83.560 128.290 83.920 131.890 ;
        RECT 84.640 131.890 86.080 133.090 ;
        RECT 84.640 128.290 85.000 131.890 ;
        RECT 85.720 128.290 86.080 131.890 ;
        RECT 86.800 131.890 88.240 133.090 ;
        RECT 86.800 128.290 87.160 131.890 ;
        RECT 87.880 128.290 88.240 131.890 ;
        RECT 88.960 131.890 90.400 133.090 ;
        RECT 88.960 128.290 89.320 131.890 ;
        RECT 90.040 128.290 90.400 131.890 ;
        RECT 91.120 131.890 92.560 133.090 ;
        RECT 91.120 128.290 91.480 131.890 ;
        RECT 92.200 128.290 92.560 131.890 ;
        RECT 93.280 131.890 94.720 133.090 ;
        RECT 93.280 128.290 93.640 131.890 ;
        RECT 94.360 128.290 94.720 131.890 ;
        RECT 95.440 131.890 96.880 133.090 ;
        RECT 95.440 128.290 95.800 131.890 ;
        RECT 96.520 128.290 96.880 131.890 ;
        RECT 97.600 131.890 99.040 133.090 ;
        RECT 97.600 128.290 97.960 131.890 ;
        RECT 100.220 124.270 102.400 133.790 ;
        RECT 111.150 133.740 111.450 134.640 ;
        RECT 113.700 134.190 114.600 135.040 ;
        RECT 118.500 140.930 151.140 153.290 ;
        RECT 153.400 151.290 153.760 154.890 ;
        RECT 154.480 154.890 155.920 156.090 ;
        RECT 154.480 151.290 154.840 154.890 ;
        RECT 155.560 151.290 155.920 154.890 ;
        RECT 156.640 154.890 158.080 156.090 ;
        RECT 156.640 151.290 157.000 154.890 ;
        RECT 153.400 141.690 154.840 144.090 ;
        RECT 155.560 141.690 157.000 144.090 ;
        RECT 159.260 140.930 160.500 156.850 ;
        RECT 118.500 139.790 160.500 140.930 ;
        RECT 118.500 136.290 146.500 139.790 ;
        RECT 106.560 132.790 107.520 133.430 ;
        RECT 118.500 132.790 127.000 136.290 ;
        RECT 103.360 131.830 104.960 132.230 ;
        RECT 102.720 130.630 103.040 131.830 ;
        RECT 104.000 131.030 105.600 131.430 ;
        RECT 105.920 130.630 106.240 131.830 ;
        RECT 103.360 130.230 104.960 130.630 ;
        RECT 103.360 127.030 104.960 127.430 ;
        RECT 102.720 125.830 103.040 127.030 ;
        RECT 104.000 126.230 105.600 126.630 ;
        RECT 105.920 125.830 106.240 127.030 ;
        RECT 103.360 125.430 104.960 125.830 ;
        RECT 106.560 124.270 127.000 132.790 ;
        RECT 100.220 121.790 127.000 124.270 ;
        RECT 81.400 118.690 82.840 121.090 ;
        RECT 83.560 118.690 85.000 121.090 ;
        RECT 85.720 118.690 87.160 121.090 ;
        RECT 87.880 118.690 89.320 121.090 ;
        RECT 90.040 118.690 91.480 121.090 ;
        RECT 92.200 118.690 93.640 121.090 ;
        RECT 94.360 118.690 95.800 121.090 ;
        RECT 96.520 118.690 97.960 121.090 ;
        RECT 100.220 117.930 101.000 121.790 ;
        RECT 54.500 117.290 101.000 117.930 ;
        RECT 74.290 96.940 75.250 102.370 ;
        RECT 76.210 100.300 78.450 100.700 ;
        RECT 75.570 98.300 75.890 99.500 ;
        RECT 76.850 98.700 79.090 99.100 ;
        RECT 79.410 98.300 79.730 99.500 ;
        RECT 76.210 97.100 78.450 97.500 ;
        RECT 80.050 96.940 81.010 102.370 ;
        RECT 91.340 102.320 121.170 102.480 ;
        RECT 74.270 96.700 75.250 96.940 ;
        RECT 80.030 96.700 81.010 96.940 ;
        RECT 90.670 101.920 121.170 102.320 ;
        RECT 90.670 101.760 99.910 101.920 ;
        RECT 63.130 91.050 64.090 95.180 ;
        RECT 65.050 94.380 67.290 94.780 ;
        RECT 64.410 92.380 64.730 93.580 ;
        RECT 65.690 92.780 67.930 93.180 ;
        RECT 68.250 92.380 68.570 93.580 ;
        RECT 65.050 91.180 67.290 91.580 ;
        RECT 68.890 91.050 69.850 95.180 ;
        RECT 74.270 92.950 75.230 96.700 ;
        RECT 76.190 96.140 78.430 96.540 ;
        RECT 75.550 94.140 75.870 95.340 ;
        RECT 76.830 94.540 79.070 94.940 ;
        RECT 79.390 94.140 79.710 95.340 ;
        RECT 74.270 92.540 75.270 92.950 ;
        RECT 76.190 92.940 78.430 93.340 ;
        RECT 80.030 92.950 80.990 96.700 ;
        RECT 63.120 90.780 64.090 91.050 ;
        RECT 68.880 90.780 69.850 91.050 ;
        RECT 63.120 87.050 64.080 90.780 ;
        RECT 65.040 90.250 67.280 90.650 ;
        RECT 64.400 88.250 64.720 89.450 ;
        RECT 65.680 88.650 67.920 89.050 ;
        RECT 68.240 88.250 68.560 89.450 ;
        RECT 65.040 87.050 67.280 87.450 ;
        RECT 68.880 87.050 69.840 90.780 ;
        RECT 74.310 88.790 75.270 92.540 ;
        RECT 76.230 92.150 78.470 92.550 ;
        RECT 80.030 92.540 81.030 92.950 ;
        RECT 75.590 90.150 75.910 91.350 ;
        RECT 76.870 90.550 79.110 90.950 ;
        RECT 79.430 90.150 79.750 91.350 ;
        RECT 76.230 88.950 78.470 89.350 ;
        RECT 80.070 88.790 81.030 92.540 ;
        RECT 74.270 88.550 75.270 88.790 ;
        RECT 80.030 88.550 81.030 88.790 ;
        RECT 63.120 86.650 64.110 87.050 ;
        RECT 68.880 86.650 69.870 87.050 ;
        RECT 63.150 82.920 64.110 86.650 ;
        RECT 65.070 86.250 67.310 86.650 ;
        RECT 64.430 84.250 64.750 85.450 ;
        RECT 65.710 84.650 67.950 85.050 ;
        RECT 68.270 84.250 68.590 85.450 ;
        RECT 65.070 83.050 67.310 83.450 ;
        RECT 68.910 82.920 69.870 86.650 ;
        RECT 74.270 84.790 75.230 88.550 ;
        RECT 76.190 87.990 78.430 88.390 ;
        RECT 75.550 85.990 75.870 87.190 ;
        RECT 76.830 86.390 79.070 86.790 ;
        RECT 79.390 85.990 79.710 87.190 ;
        RECT 76.190 84.790 78.430 85.190 ;
        RECT 80.030 84.790 80.990 88.550 ;
        RECT 90.670 85.840 91.230 101.760 ;
        RECT 91.790 99.800 93.850 101.000 ;
        RECT 93.490 96.200 93.850 99.800 ;
        RECT 94.570 99.800 96.010 101.000 ;
        RECT 94.570 96.200 94.930 99.800 ;
        RECT 95.650 96.200 96.010 99.800 ;
        RECT 96.730 99.800 98.700 101.000 ;
        RECT 96.730 96.200 97.090 99.800 ;
        RECT 93.490 86.600 94.930 89.000 ;
        RECT 95.650 86.600 97.090 89.000 ;
        RECT 99.350 85.840 99.910 101.760 ;
        RECT 90.670 85.490 99.910 85.840 ;
        RECT 101.340 101.840 110.580 101.920 ;
        RECT 101.340 85.920 101.900 101.840 ;
        RECT 102.440 99.880 104.520 101.080 ;
        RECT 104.160 96.280 104.520 99.880 ;
        RECT 105.240 99.880 106.680 101.080 ;
        RECT 105.240 96.280 105.600 99.880 ;
        RECT 106.320 96.280 106.680 99.880 ;
        RECT 107.400 99.880 109.480 101.080 ;
        RECT 107.400 96.280 107.760 99.880 ;
        RECT 104.160 86.680 105.600 89.080 ;
        RECT 106.320 86.680 107.760 89.080 ;
        RECT 110.020 85.920 110.580 101.840 ;
        RECT 101.340 85.490 110.580 85.920 ;
        RECT 111.930 86.000 112.490 101.920 ;
        RECT 118.170 101.160 119.370 101.920 ;
        RECT 113.060 99.960 115.110 101.160 ;
        RECT 114.750 96.360 115.110 99.960 ;
        RECT 115.830 99.960 117.270 101.160 ;
        RECT 115.830 96.360 116.190 99.960 ;
        RECT 116.910 96.360 117.270 99.960 ;
        RECT 117.990 99.960 120.100 101.160 ;
        RECT 117.990 96.360 118.350 99.960 ;
        RECT 114.750 86.760 116.190 89.160 ;
        RECT 116.910 86.760 118.350 89.160 ;
        RECT 120.610 86.000 121.170 101.920 ;
        RECT 111.930 85.490 121.170 86.000 ;
        RECT 90.670 85.280 159.450 85.490 ;
        RECT 74.270 84.390 75.250 84.790 ;
        RECT 80.030 84.390 81.010 84.790 ;
        RECT 63.140 82.650 64.110 82.920 ;
        RECT 68.900 82.650 69.870 82.920 ;
        RECT 63.140 78.930 64.100 82.650 ;
        RECT 65.060 82.120 67.300 82.520 ;
        RECT 64.420 80.120 64.740 81.320 ;
        RECT 65.700 80.520 67.940 80.920 ;
        RECT 68.260 80.120 68.580 81.320 ;
        RECT 63.140 78.520 64.110 78.930 ;
        RECT 65.060 78.920 67.300 79.320 ;
        RECT 68.900 78.930 69.860 82.650 ;
        RECT 74.290 80.630 75.250 84.390 ;
        RECT 76.210 83.990 78.450 84.390 ;
        RECT 75.570 81.990 75.890 83.190 ;
        RECT 76.850 82.390 79.090 82.790 ;
        RECT 79.410 81.990 79.730 83.190 ;
        RECT 76.210 80.790 78.450 81.190 ;
        RECT 80.050 80.630 81.010 84.390 ;
        RECT 74.270 80.390 75.250 80.630 ;
        RECT 80.030 80.390 81.010 80.630 ;
        RECT 63.150 74.800 64.110 78.520 ;
        RECT 65.070 78.130 67.310 78.530 ;
        RECT 68.900 78.520 69.870 78.930 ;
        RECT 64.430 76.130 64.750 77.330 ;
        RECT 65.710 76.530 67.950 76.930 ;
        RECT 68.270 76.130 68.590 77.330 ;
        RECT 65.070 74.930 67.310 75.330 ;
        RECT 68.910 74.800 69.870 78.520 ;
        RECT 74.270 76.500 75.230 80.390 ;
        RECT 76.190 79.830 78.430 80.230 ;
        RECT 75.550 77.830 75.870 79.030 ;
        RECT 76.830 78.230 79.070 78.630 ;
        RECT 79.390 77.830 79.710 79.030 ;
        RECT 76.190 76.630 78.430 77.030 ;
        RECT 80.030 76.500 80.990 80.390 ;
        RECT 90.800 77.390 159.450 85.280 ;
        RECT 92.690 76.920 159.450 77.390 ;
        RECT 74.270 76.230 75.250 76.500 ;
        RECT 80.030 76.230 81.010 76.500 ;
        RECT 63.140 74.530 64.110 74.800 ;
        RECT 68.900 74.530 69.870 74.800 ;
        RECT 35.810 73.640 36.770 73.660 ;
        RECT 4.760 73.440 26.960 73.550 ;
        RECT 33.890 73.540 40.640 73.640 ;
        RECT 0.580 72.990 26.960 73.440 ;
        RECT 0.580 57.070 5.410 72.990 ;
        RECT 6.500 71.030 7.940 72.230 ;
        RECT 7.580 67.430 7.940 71.030 ;
        RECT 8.660 71.030 10.100 72.230 ;
        RECT 8.660 67.430 9.020 71.030 ;
        RECT 9.740 67.430 10.100 71.030 ;
        RECT 10.820 71.030 12.260 72.230 ;
        RECT 10.820 67.430 11.180 71.030 ;
        RECT 11.900 67.430 12.260 71.030 ;
        RECT 12.980 71.030 14.420 72.230 ;
        RECT 12.980 67.430 13.340 71.030 ;
        RECT 14.060 67.430 14.420 71.030 ;
        RECT 15.140 71.030 16.580 72.230 ;
        RECT 15.140 67.430 15.500 71.030 ;
        RECT 16.220 67.430 16.580 71.030 ;
        RECT 17.300 71.030 18.740 72.230 ;
        RECT 17.300 67.430 17.660 71.030 ;
        RECT 18.380 67.430 18.740 71.030 ;
        RECT 19.460 71.030 20.900 72.230 ;
        RECT 19.460 67.430 19.820 71.030 ;
        RECT 20.540 67.430 20.900 71.030 ;
        RECT 21.620 71.030 23.060 72.230 ;
        RECT 21.620 67.430 21.980 71.030 ;
        RECT 22.700 67.430 23.060 71.030 ;
        RECT 23.780 71.030 25.220 72.230 ;
        RECT 23.780 67.430 24.140 71.030 ;
        RECT 7.580 57.830 9.020 60.230 ;
        RECT 9.740 57.830 11.180 60.230 ;
        RECT 11.900 57.830 13.340 60.230 ;
        RECT 14.060 57.830 15.500 60.230 ;
        RECT 16.220 57.830 17.660 60.230 ;
        RECT 18.380 57.830 19.820 60.230 ;
        RECT 20.540 57.830 21.980 60.230 ;
        RECT 22.700 57.830 24.140 60.230 ;
        RECT 26.400 57.070 26.960 72.990 ;
        RECT 33.880 72.680 40.640 73.540 ;
        RECT 33.880 72.580 40.610 72.680 ;
        RECT 33.890 69.540 34.850 72.580 ;
        RECT 35.810 69.680 36.770 72.580 ;
        RECT 39.650 69.540 40.610 72.580 ;
        RECT 63.140 70.790 64.100 74.530 ;
        RECT 65.060 74.000 67.300 74.400 ;
        RECT 64.420 72.000 64.740 73.200 ;
        RECT 65.700 72.400 67.940 72.800 ;
        RECT 68.260 72.000 68.580 73.200 ;
        RECT 65.060 70.800 67.300 71.200 ;
        RECT 68.900 70.790 69.860 74.530 ;
        RECT 74.290 72.340 75.250 76.230 ;
        RECT 76.210 75.700 78.450 76.100 ;
        RECT 75.570 73.700 75.890 74.900 ;
        RECT 76.850 74.100 79.090 74.500 ;
        RECT 79.410 73.700 79.730 74.900 ;
        RECT 76.210 72.500 78.450 72.900 ;
        RECT 80.050 72.340 81.010 76.230 ;
        RECT 74.290 72.100 75.260 72.340 ;
        RECT 80.050 72.100 81.020 72.340 ;
        RECT 63.140 70.400 64.130 70.790 ;
        RECT 68.900 70.400 69.890 70.790 ;
        RECT 33.880 68.390 34.850 69.540 ;
        RECT 35.800 68.740 38.040 69.140 ;
        RECT 33.880 65.630 34.840 68.390 ;
        RECT 39.640 68.160 40.610 69.540 ;
        RECT 35.160 66.740 35.480 67.940 ;
        RECT 36.440 67.140 38.680 67.540 ;
        RECT 39.000 66.740 39.320 67.940 ;
        RECT 33.880 65.140 34.870 65.630 ;
        RECT 35.800 65.540 38.040 65.940 ;
        RECT 39.640 65.910 40.600 68.160 ;
        RECT 63.170 66.660 64.130 70.400 ;
        RECT 65.090 69.990 67.330 70.390 ;
        RECT 64.450 67.990 64.770 69.190 ;
        RECT 65.730 68.390 67.970 68.790 ;
        RECT 68.290 67.990 68.610 69.190 ;
        RECT 65.090 66.790 67.330 67.190 ;
        RECT 68.930 66.660 69.890 70.400 ;
        RECT 74.300 68.210 75.260 72.100 ;
        RECT 76.220 71.540 78.460 71.940 ;
        RECT 75.580 69.540 75.900 70.740 ;
        RECT 76.860 69.940 79.100 70.340 ;
        RECT 79.420 69.540 79.740 70.740 ;
        RECT 76.220 68.340 78.460 68.740 ;
        RECT 80.060 68.210 81.020 72.100 ;
        RECT 63.160 66.390 64.130 66.660 ;
        RECT 68.920 66.390 69.890 66.660 ;
        RECT 74.280 67.940 75.260 68.210 ;
        RECT 80.040 67.940 81.020 68.210 ;
        RECT 39.640 65.140 40.630 65.910 ;
        RECT 33.910 64.520 34.870 65.140 ;
        RECT 39.670 64.520 40.630 65.140 ;
        RECT 33.900 62.790 34.870 64.520 ;
        RECT 35.820 63.720 38.060 64.120 ;
        RECT 33.900 60.120 34.860 62.790 ;
        RECT 35.180 61.720 35.500 62.920 ;
        RECT 36.460 62.120 38.700 62.520 ;
        RECT 39.020 61.720 39.340 62.920 ;
        RECT 39.660 62.810 40.630 64.520 ;
        RECT 35.820 60.520 38.060 60.920 ;
        RECT 39.660 60.120 40.620 62.810 ;
        RECT 63.160 62.670 64.120 66.390 ;
        RECT 65.080 65.860 67.320 66.260 ;
        RECT 64.440 63.860 64.760 65.060 ;
        RECT 65.720 64.260 67.960 64.660 ;
        RECT 68.280 63.860 68.600 65.060 ;
        RECT 63.160 62.260 64.130 62.670 ;
        RECT 65.080 62.660 67.320 63.060 ;
        RECT 68.920 62.670 69.880 66.390 ;
        RECT 74.280 64.050 75.240 67.940 ;
        RECT 76.200 67.410 78.440 67.810 ;
        RECT 75.560 65.410 75.880 66.610 ;
        RECT 76.840 65.810 79.080 66.210 ;
        RECT 79.400 65.410 79.720 66.610 ;
        RECT 76.200 64.210 78.440 64.610 ;
        RECT 80.040 64.050 81.000 67.940 ;
        RECT 74.280 63.810 75.260 64.050 ;
        RECT 80.040 63.810 81.020 64.050 ;
        RECT 0.580 56.510 26.960 57.070 ;
        RECT 0.580 55.960 5.410 56.510 ;
        RECT 0.580 55.400 26.860 55.960 ;
        RECT 0.580 39.480 5.410 55.400 ;
        RECT 6.400 53.440 7.840 54.640 ;
        RECT 7.480 49.840 7.840 53.440 ;
        RECT 8.560 53.440 10.000 54.640 ;
        RECT 8.560 49.840 8.920 53.440 ;
        RECT 9.640 49.840 10.000 53.440 ;
        RECT 10.720 53.440 12.160 54.640 ;
        RECT 10.720 49.840 11.080 53.440 ;
        RECT 11.800 49.840 12.160 53.440 ;
        RECT 12.880 53.440 14.320 54.640 ;
        RECT 12.880 49.840 13.240 53.440 ;
        RECT 13.960 49.840 14.320 53.440 ;
        RECT 15.040 53.440 16.480 54.640 ;
        RECT 15.040 49.840 15.400 53.440 ;
        RECT 16.120 49.840 16.480 53.440 ;
        RECT 17.200 53.440 18.640 54.640 ;
        RECT 17.200 49.840 17.560 53.440 ;
        RECT 18.280 49.840 18.640 53.440 ;
        RECT 19.360 53.440 20.800 54.640 ;
        RECT 19.360 49.840 19.720 53.440 ;
        RECT 20.440 49.840 20.800 53.440 ;
        RECT 21.520 53.440 22.960 54.640 ;
        RECT 21.520 49.840 21.880 53.440 ;
        RECT 22.600 49.840 22.960 53.440 ;
        RECT 23.680 53.440 25.120 54.640 ;
        RECT 23.680 49.840 24.040 53.440 ;
        RECT 7.480 40.240 8.920 42.640 ;
        RECT 9.640 40.240 11.080 42.640 ;
        RECT 11.800 40.240 13.240 42.640 ;
        RECT 13.960 40.240 15.400 42.640 ;
        RECT 16.120 40.240 17.560 42.640 ;
        RECT 18.280 40.240 19.720 42.640 ;
        RECT 20.440 40.240 21.880 42.640 ;
        RECT 22.600 40.240 24.040 42.640 ;
        RECT 26.300 39.480 26.860 55.400 ;
        RECT 29.130 49.170 30.090 58.940 ;
        RECT 31.050 56.670 33.290 57.070 ;
        RECT 30.410 54.670 30.730 55.870 ;
        RECT 31.690 55.070 33.930 55.470 ;
        RECT 34.250 54.670 34.570 55.870 ;
        RECT 31.050 53.470 33.290 53.870 ;
        RECT 31.050 52.560 33.290 52.960 ;
        RECT 30.410 50.560 30.730 51.760 ;
        RECT 31.690 50.960 33.930 51.360 ;
        RECT 34.250 50.560 34.570 51.760 ;
        RECT 31.050 49.360 33.290 49.760 ;
        RECT 34.890 49.170 35.850 58.870 ;
        RECT 39.040 49.210 40.000 58.870 ;
        RECT 40.960 56.710 43.200 57.110 ;
        RECT 40.320 54.710 40.640 55.910 ;
        RECT 41.600 55.110 43.840 55.510 ;
        RECT 44.160 54.710 44.480 55.910 ;
        RECT 40.960 53.510 43.200 53.910 ;
        RECT 40.960 52.600 43.200 53.000 ;
        RECT 40.320 50.600 40.640 51.800 ;
        RECT 41.600 51.000 43.840 51.400 ;
        RECT 44.160 50.600 44.480 51.800 ;
        RECT 40.960 49.400 43.200 49.800 ;
        RECT 44.800 49.210 45.760 58.940 ;
        RECT 54.660 54.830 55.620 61.000 ;
        RECT 56.580 58.430 58.820 58.830 ;
        RECT 55.940 56.430 56.260 57.630 ;
        RECT 57.220 56.830 59.460 57.230 ;
        RECT 59.780 56.430 60.100 57.630 ;
        RECT 56.580 55.230 58.820 55.630 ;
        RECT 60.420 54.830 61.380 61.060 ;
        RECT 63.170 58.540 64.130 62.260 ;
        RECT 65.090 61.870 67.330 62.270 ;
        RECT 68.920 62.260 69.890 62.670 ;
        RECT 64.450 59.870 64.770 61.070 ;
        RECT 65.730 60.270 67.970 60.670 ;
        RECT 68.290 59.870 68.610 61.070 ;
        RECT 65.090 58.670 67.330 59.070 ;
        RECT 68.930 58.540 69.890 62.260 ;
        RECT 74.300 59.650 75.260 63.810 ;
        RECT 76.220 63.250 78.460 63.650 ;
        RECT 75.580 61.250 75.900 62.450 ;
        RECT 76.860 61.650 79.100 62.050 ;
        RECT 79.420 61.250 79.740 62.450 ;
        RECT 76.220 60.050 78.460 60.450 ;
        RECT 80.060 59.650 81.020 63.810 ;
        RECT 83.650 59.650 84.610 65.790 ;
        RECT 85.570 63.250 87.810 63.650 ;
        RECT 84.930 61.250 85.250 62.450 ;
        RECT 86.210 61.650 88.450 62.050 ;
        RECT 88.770 61.250 89.090 62.450 ;
        RECT 85.570 60.050 87.810 60.450 ;
        RECT 89.410 59.650 90.370 65.760 ;
        RECT 63.160 58.270 64.130 58.540 ;
        RECT 68.920 58.270 69.890 58.540 ;
        RECT 29.120 48.960 30.090 49.170 ;
        RECT 34.880 48.960 35.850 49.170 ;
        RECT 39.030 49.000 40.000 49.210 ;
        RECT 44.790 49.000 45.760 49.210 ;
        RECT 54.910 53.380 59.410 53.420 ;
        RECT 63.160 53.380 64.120 58.270 ;
        RECT 65.080 57.740 67.320 58.140 ;
        RECT 64.440 55.740 64.760 56.940 ;
        RECT 65.720 56.140 67.960 56.540 ;
        RECT 68.280 55.740 68.600 56.940 ;
        RECT 65.080 54.540 67.320 54.940 ;
        RECT 68.920 53.430 69.880 58.270 ;
        RECT 74.230 53.430 75.190 58.530 ;
        RECT 76.150 57.730 78.390 58.130 ;
        RECT 75.510 55.730 75.830 56.930 ;
        RECT 76.790 56.130 79.030 56.530 ;
        RECT 79.350 55.730 79.670 56.930 ;
        RECT 76.150 54.530 78.390 54.930 ;
        RECT 76.150 53.430 77.110 53.980 ;
        RECT 79.990 53.430 80.950 58.530 ;
        RECT 65.040 53.380 80.950 53.430 ;
        RECT 54.910 52.630 80.950 53.380 ;
        RECT 54.910 51.130 81.300 52.630 ;
        RECT 92.690 51.130 93.890 76.920 ;
        RECT 149.920 76.910 159.450 76.920 ;
        RECT 138.520 72.440 139.580 74.520 ;
        RECT 138.490 71.280 139.580 72.440 ;
        RECT 138.490 70.120 139.550 71.280 ;
        RECT 138.160 70.100 139.550 70.120 ;
        RECT 107.110 69.690 129.310 70.010 ;
        RECT 136.240 70.000 142.990 70.100 ;
        RECT 105.580 69.450 129.310 69.690 ;
        RECT 105.580 53.530 107.670 69.450 ;
        RECT 108.850 67.490 110.290 68.690 ;
        RECT 109.930 63.890 110.290 67.490 ;
        RECT 111.010 67.490 112.450 68.690 ;
        RECT 111.010 63.890 111.370 67.490 ;
        RECT 112.090 63.890 112.450 67.490 ;
        RECT 113.170 67.490 114.610 68.690 ;
        RECT 113.170 63.890 113.530 67.490 ;
        RECT 114.250 63.890 114.610 67.490 ;
        RECT 115.330 67.490 116.770 68.690 ;
        RECT 115.330 63.890 115.690 67.490 ;
        RECT 116.410 63.890 116.770 67.490 ;
        RECT 117.490 67.490 118.930 68.690 ;
        RECT 117.490 63.890 117.850 67.490 ;
        RECT 118.570 63.890 118.930 67.490 ;
        RECT 119.650 67.490 121.090 68.690 ;
        RECT 119.650 63.890 120.010 67.490 ;
        RECT 120.730 63.890 121.090 67.490 ;
        RECT 121.810 67.490 123.250 68.690 ;
        RECT 121.810 63.890 122.170 67.490 ;
        RECT 122.890 63.890 123.250 67.490 ;
        RECT 123.970 67.490 125.410 68.690 ;
        RECT 123.970 63.890 124.330 67.490 ;
        RECT 125.050 63.890 125.410 67.490 ;
        RECT 126.130 67.490 127.570 68.690 ;
        RECT 126.130 63.890 126.490 67.490 ;
        RECT 109.930 54.290 111.370 56.690 ;
        RECT 112.090 54.290 113.530 56.690 ;
        RECT 114.250 54.290 115.690 56.690 ;
        RECT 116.410 54.290 117.850 56.690 ;
        RECT 118.570 54.290 120.010 56.690 ;
        RECT 120.730 54.290 122.170 56.690 ;
        RECT 122.890 54.290 124.330 56.690 ;
        RECT 125.050 54.290 126.490 56.690 ;
        RECT 128.750 53.530 129.310 69.450 ;
        RECT 136.230 69.140 142.990 70.000 ;
        RECT 136.230 69.040 142.960 69.140 ;
        RECT 136.240 66.000 137.200 69.040 ;
        RECT 138.160 66.140 139.120 69.040 ;
        RECT 142.000 66.000 142.960 69.040 ;
        RECT 136.230 64.850 137.200 66.000 ;
        RECT 138.150 65.200 140.390 65.600 ;
        RECT 136.230 62.090 137.190 64.850 ;
        RECT 141.990 64.620 142.960 66.000 ;
        RECT 137.510 63.200 137.830 64.400 ;
        RECT 138.790 63.600 141.030 64.000 ;
        RECT 141.350 63.200 141.670 64.400 ;
        RECT 136.230 61.600 137.220 62.090 ;
        RECT 138.150 62.000 140.390 62.400 ;
        RECT 141.990 62.370 142.950 64.620 ;
        RECT 141.990 61.600 142.980 62.370 ;
        RECT 136.260 60.980 137.220 61.600 ;
        RECT 142.020 60.980 142.980 61.600 ;
        RECT 136.250 59.250 137.220 60.980 ;
        RECT 138.170 60.180 140.410 60.580 ;
        RECT 136.250 56.580 137.210 59.250 ;
        RECT 137.530 58.180 137.850 59.380 ;
        RECT 138.810 58.580 141.050 58.980 ;
        RECT 141.370 58.180 141.690 59.380 ;
        RECT 142.010 59.270 142.980 60.980 ;
        RECT 138.170 56.980 140.410 57.380 ;
        RECT 142.010 56.580 142.970 59.270 ;
        RECT 105.580 52.970 129.310 53.530 ;
        RECT 105.580 52.420 107.670 52.970 ;
        RECT 105.580 51.860 129.210 52.420 ;
        RECT 105.580 51.850 107.670 51.860 ;
        RECT 54.910 50.570 94.190 51.130 ;
        RECT 54.910 50.550 81.300 50.570 ;
        RECT 29.120 40.660 30.080 48.960 ;
        RECT 31.040 48.370 33.280 48.770 ;
        RECT 30.400 46.370 30.720 47.570 ;
        RECT 31.680 46.770 33.920 47.170 ;
        RECT 34.240 46.370 34.560 47.570 ;
        RECT 31.040 45.170 33.280 45.570 ;
        RECT 31.040 44.260 33.280 44.660 ;
        RECT 30.400 42.260 30.720 43.460 ;
        RECT 31.680 42.660 33.920 43.060 ;
        RECT 34.240 42.260 34.560 43.460 ;
        RECT 31.040 41.060 33.280 41.460 ;
        RECT 34.880 40.660 35.840 48.960 ;
        RECT 39.030 40.700 39.990 49.000 ;
        RECT 40.950 48.410 43.190 48.810 ;
        RECT 40.310 46.410 40.630 47.610 ;
        RECT 41.590 46.810 43.830 47.210 ;
        RECT 44.150 46.410 44.470 47.610 ;
        RECT 40.950 45.210 43.190 45.610 ;
        RECT 40.950 44.300 43.190 44.700 ;
        RECT 40.310 42.300 40.630 43.500 ;
        RECT 41.590 42.700 43.830 43.100 ;
        RECT 44.150 42.300 44.470 43.500 ;
        RECT 40.950 41.100 43.190 41.500 ;
        RECT 44.790 40.700 45.750 49.000 ;
        RECT 0.580 38.920 26.860 39.480 ;
        RECT 0.580 38.490 5.410 38.920 ;
        RECT 0.580 37.930 26.800 38.490 ;
        RECT 0.580 22.010 5.410 37.930 ;
        RECT 6.340 35.970 7.780 37.170 ;
        RECT 7.420 32.370 7.780 35.970 ;
        RECT 8.500 35.970 9.940 37.170 ;
        RECT 8.500 32.370 8.860 35.970 ;
        RECT 9.580 32.370 9.940 35.970 ;
        RECT 10.660 35.970 12.100 37.170 ;
        RECT 10.660 32.370 11.020 35.970 ;
        RECT 11.740 32.370 12.100 35.970 ;
        RECT 12.820 35.970 14.260 37.170 ;
        RECT 12.820 32.370 13.180 35.970 ;
        RECT 13.900 32.370 14.260 35.970 ;
        RECT 14.980 35.970 16.420 37.170 ;
        RECT 14.980 32.370 15.340 35.970 ;
        RECT 16.060 32.370 16.420 35.970 ;
        RECT 17.140 35.970 18.580 37.170 ;
        RECT 17.140 32.370 17.500 35.970 ;
        RECT 18.220 32.370 18.580 35.970 ;
        RECT 19.300 35.970 20.740 37.170 ;
        RECT 19.300 32.370 19.660 35.970 ;
        RECT 20.380 32.370 20.740 35.970 ;
        RECT 21.460 35.970 22.900 37.170 ;
        RECT 21.460 32.370 21.820 35.970 ;
        RECT 22.540 32.370 22.900 35.970 ;
        RECT 23.620 35.970 25.060 37.170 ;
        RECT 23.620 32.370 23.980 35.970 ;
        RECT 7.420 22.770 8.860 25.170 ;
        RECT 9.580 22.770 11.020 25.170 ;
        RECT 11.740 22.770 13.180 25.170 ;
        RECT 13.900 22.770 15.340 25.170 ;
        RECT 16.060 22.770 17.500 25.170 ;
        RECT 18.220 22.770 19.660 25.170 ;
        RECT 20.380 22.770 21.820 25.170 ;
        RECT 22.540 22.770 23.980 25.170 ;
        RECT 26.240 22.010 26.800 37.930 ;
        RECT 29.130 30.310 30.090 37.300 ;
        RECT 31.050 36.500 33.290 36.900 ;
        RECT 30.410 34.500 30.730 35.700 ;
        RECT 31.690 34.900 33.930 35.300 ;
        RECT 34.250 34.500 34.570 35.700 ;
        RECT 31.050 33.300 33.290 33.700 ;
        RECT 31.050 30.310 32.010 32.190 ;
        RECT 34.890 30.310 35.850 37.300 ;
        RECT 39.050 30.310 40.010 37.290 ;
        RECT 40.970 36.490 43.210 36.890 ;
        RECT 40.330 34.490 40.650 35.690 ;
        RECT 41.610 34.890 43.850 35.290 ;
        RECT 44.170 34.490 44.490 35.690 ;
        RECT 40.970 33.290 43.210 33.690 ;
        RECT 40.970 30.310 41.930 32.310 ;
        RECT 44.810 30.310 45.770 37.290 ;
        RECT 29.130 30.300 45.770 30.310 ;
        RECT 0.580 21.600 26.800 22.010 ;
        RECT 28.970 29.330 45.770 30.300 ;
        RECT 54.910 33.480 59.410 50.550 ;
        RECT 66.070 45.950 67.030 46.000 ;
        RECT 62.250 44.990 67.030 45.950 ;
        RECT 60.310 39.500 61.270 44.760 ;
        RECT 62.230 42.820 64.470 43.220 ;
        RECT 61.590 40.820 61.910 42.020 ;
        RECT 62.870 41.220 65.110 41.620 ;
        RECT 65.430 40.820 65.750 42.020 ;
        RECT 62.230 39.620 64.470 40.020 ;
        RECT 66.070 39.500 67.030 44.990 ;
        RECT 60.310 39.220 61.280 39.500 ;
        RECT 66.070 39.220 67.040 39.500 ;
        RECT 60.320 35.100 61.280 39.220 ;
        RECT 62.240 38.700 64.480 39.100 ;
        RECT 61.600 36.700 61.920 37.900 ;
        RECT 62.880 37.100 65.120 37.500 ;
        RECT 65.440 36.700 65.760 37.900 ;
        RECT 62.240 35.500 64.480 35.900 ;
        RECT 66.080 35.100 67.040 39.220 ;
        RECT 70.860 34.730 71.420 50.550 ;
        RECT 71.930 48.690 74.040 49.890 ;
        RECT 73.680 45.090 74.040 48.690 ;
        RECT 74.760 48.690 76.200 49.890 ;
        RECT 74.760 45.090 75.120 48.690 ;
        RECT 75.840 45.090 76.200 48.690 ;
        RECT 76.920 48.690 79.000 49.890 ;
        RECT 76.920 45.090 77.280 48.690 ;
        RECT 73.680 35.490 75.120 37.890 ;
        RECT 75.840 35.490 77.280 37.890 ;
        RECT 79.540 34.730 80.100 50.550 ;
        RECT 70.860 34.410 80.100 34.730 ;
        RECT 80.630 34.650 81.190 50.550 ;
        RECT 81.650 49.810 83.520 49.880 ;
        RECT 81.650 48.680 83.810 49.810 ;
        RECT 82.370 48.610 83.810 48.680 ;
        RECT 83.450 45.010 83.810 48.610 ;
        RECT 84.530 48.610 85.970 49.810 ;
        RECT 84.530 45.010 84.890 48.610 ;
        RECT 85.610 45.010 85.970 48.610 ;
        RECT 86.690 48.610 88.130 49.810 ;
        RECT 86.690 45.010 87.050 48.610 ;
        RECT 87.770 45.010 88.130 48.610 ;
        RECT 88.850 48.610 90.290 49.810 ;
        RECT 88.850 45.010 89.210 48.610 ;
        RECT 89.930 45.010 90.290 48.610 ;
        RECT 91.010 48.610 92.960 49.810 ;
        RECT 91.010 45.010 91.370 48.610 ;
        RECT 83.450 35.410 84.890 37.810 ;
        RECT 85.610 35.410 87.050 37.810 ;
        RECT 87.770 35.410 89.210 37.810 ;
        RECT 89.930 35.410 91.370 37.810 ;
        RECT 93.630 34.650 94.190 50.570 ;
        RECT 80.630 34.410 94.190 34.650 ;
        RECT 105.580 35.940 107.570 51.850 ;
        RECT 108.750 49.900 110.190 51.100 ;
        RECT 109.830 46.300 110.190 49.900 ;
        RECT 110.910 49.900 112.350 51.100 ;
        RECT 110.910 46.300 111.270 49.900 ;
        RECT 111.990 46.300 112.350 49.900 ;
        RECT 113.070 49.900 114.510 51.100 ;
        RECT 113.070 46.300 113.430 49.900 ;
        RECT 114.150 46.300 114.510 49.900 ;
        RECT 115.230 49.900 116.670 51.100 ;
        RECT 115.230 46.300 115.590 49.900 ;
        RECT 116.310 46.300 116.670 49.900 ;
        RECT 117.390 49.900 118.830 51.100 ;
        RECT 117.390 46.300 117.750 49.900 ;
        RECT 118.470 46.300 118.830 49.900 ;
        RECT 119.550 49.900 120.990 51.100 ;
        RECT 119.550 46.300 119.910 49.900 ;
        RECT 120.630 46.300 120.990 49.900 ;
        RECT 121.710 49.900 123.150 51.100 ;
        RECT 121.710 46.300 122.070 49.900 ;
        RECT 122.790 46.300 123.150 49.900 ;
        RECT 123.870 49.900 125.310 51.100 ;
        RECT 123.870 46.300 124.230 49.900 ;
        RECT 124.950 46.300 125.310 49.900 ;
        RECT 126.030 49.900 127.470 51.100 ;
        RECT 126.030 46.300 126.390 49.900 ;
        RECT 109.830 36.700 111.270 39.100 ;
        RECT 111.990 36.700 113.430 39.100 ;
        RECT 114.150 36.700 115.590 39.100 ;
        RECT 116.310 36.700 117.750 39.100 ;
        RECT 118.470 36.700 119.910 39.100 ;
        RECT 120.630 36.700 122.070 39.100 ;
        RECT 122.790 36.700 124.230 39.100 ;
        RECT 124.950 36.700 126.390 39.100 ;
        RECT 128.650 35.940 129.210 51.860 ;
        RECT 131.480 45.630 132.440 55.400 ;
        RECT 133.400 53.130 135.640 53.530 ;
        RECT 132.760 51.130 133.080 52.330 ;
        RECT 134.040 51.530 136.280 51.930 ;
        RECT 136.600 51.130 136.920 52.330 ;
        RECT 133.400 49.930 135.640 50.330 ;
        RECT 133.400 49.020 135.640 49.420 ;
        RECT 132.760 47.020 133.080 48.220 ;
        RECT 134.040 47.420 136.280 47.820 ;
        RECT 136.600 47.020 136.920 48.220 ;
        RECT 133.400 45.820 135.640 46.220 ;
        RECT 137.240 45.630 138.200 55.330 ;
        RECT 141.390 45.670 142.350 55.330 ;
        RECT 143.310 53.170 145.550 53.570 ;
        RECT 142.670 51.170 142.990 52.370 ;
        RECT 143.950 51.570 146.190 51.970 ;
        RECT 146.510 51.170 146.830 52.370 ;
        RECT 143.310 49.970 145.550 50.370 ;
        RECT 143.310 49.060 145.550 49.460 ;
        RECT 142.670 47.060 142.990 48.260 ;
        RECT 143.950 47.460 146.190 47.860 ;
        RECT 146.510 47.060 146.830 48.260 ;
        RECT 143.310 45.860 145.550 46.260 ;
        RECT 147.150 45.670 148.110 55.400 ;
        RECT 131.470 45.420 132.440 45.630 ;
        RECT 137.230 45.420 138.200 45.630 ;
        RECT 141.380 45.460 142.350 45.670 ;
        RECT 147.140 45.460 148.110 45.670 ;
        RECT 131.470 37.120 132.430 45.420 ;
        RECT 133.390 44.830 135.630 45.230 ;
        RECT 132.750 42.830 133.070 44.030 ;
        RECT 134.030 43.230 136.270 43.630 ;
        RECT 136.590 42.830 136.910 44.030 ;
        RECT 133.390 41.630 135.630 42.030 ;
        RECT 133.390 40.720 135.630 41.120 ;
        RECT 132.750 38.720 133.070 39.920 ;
        RECT 134.030 39.120 136.270 39.520 ;
        RECT 136.590 38.720 136.910 39.920 ;
        RECT 133.390 37.520 135.630 37.920 ;
        RECT 137.230 37.120 138.190 45.420 ;
        RECT 141.380 37.160 142.340 45.460 ;
        RECT 143.300 44.870 145.540 45.270 ;
        RECT 142.660 42.870 142.980 44.070 ;
        RECT 143.940 43.270 146.180 43.670 ;
        RECT 146.500 42.870 146.820 44.070 ;
        RECT 143.300 41.670 145.540 42.070 ;
        RECT 143.300 40.760 145.540 41.160 ;
        RECT 142.660 38.760 142.980 39.960 ;
        RECT 143.940 39.160 146.180 39.560 ;
        RECT 146.500 38.760 146.820 39.960 ;
        RECT 143.300 37.560 145.540 37.960 ;
        RECT 147.140 37.160 148.100 45.460 ;
        RECT 105.580 35.380 129.210 35.940 ;
        RECT 105.580 34.950 107.570 35.380 ;
        RECT 62.310 33.480 64.420 33.700 ;
        RECT 69.930 33.480 94.270 34.410 ;
        RECT 54.910 32.790 94.270 33.480 ;
        RECT 105.580 34.390 129.150 34.950 ;
        RECT 54.910 31.780 71.370 32.790 ;
        RECT 28.970 24.880 45.320 29.330 ;
        RECT 54.910 25.100 59.410 31.780 ;
        RECT 62.310 25.100 64.420 31.780 ;
        RECT 68.300 29.955 74.740 30.450 ;
        RECT 68.300 25.100 68.795 29.955 ;
        RECT 69.115 29.275 73.925 29.635 ;
        RECT 69.115 25.185 69.475 29.275 ;
        RECT 69.785 25.495 73.255 28.965 ;
        RECT 73.565 25.185 73.925 29.275 ;
        RECT 69.115 25.100 73.925 25.185 ;
        RECT 74.245 25.100 74.740 29.955 ;
        RECT 76.270 29.955 82.710 30.450 ;
        RECT 76.270 25.100 76.765 29.955 ;
        RECT 77.085 29.275 81.895 29.635 ;
        RECT 77.085 25.185 77.445 29.275 ;
        RECT 77.755 25.495 81.225 28.965 ;
        RECT 81.535 25.185 81.895 29.275 ;
        RECT 77.085 25.100 81.895 25.185 ;
        RECT 82.215 25.100 82.710 29.955 ;
        RECT 84.240 29.955 90.680 30.450 ;
        RECT 84.240 25.100 84.735 29.955 ;
        RECT 85.055 29.275 89.865 29.635 ;
        RECT 85.055 25.185 85.415 29.275 ;
        RECT 85.725 25.495 89.195 28.965 ;
        RECT 89.505 25.185 89.865 29.275 ;
        RECT 85.055 25.100 89.865 25.185 ;
        RECT 90.185 25.100 90.680 29.955 ;
        RECT 54.910 24.880 90.680 25.100 ;
        RECT 28.970 24.010 90.680 24.880 ;
        RECT 28.970 21.600 64.420 24.010 ;
        RECT 0.580 17.010 64.420 21.600 ;
        RECT 68.300 21.855 74.740 22.350 ;
        RECT 68.300 17.010 68.795 21.855 ;
        RECT 69.115 21.175 73.925 21.535 ;
        RECT 69.115 17.085 69.475 21.175 ;
        RECT 69.785 17.395 73.255 20.865 ;
        RECT 73.565 17.085 73.925 21.175 ;
        RECT 69.115 17.010 73.925 17.085 ;
        RECT 74.245 17.010 74.740 21.855 ;
        RECT 76.270 21.855 82.710 22.350 ;
        RECT 76.270 17.010 76.765 21.855 ;
        RECT 77.085 21.175 81.895 21.535 ;
        RECT 77.085 17.085 77.445 21.175 ;
        RECT 77.755 17.395 81.225 20.865 ;
        RECT 81.535 17.085 81.895 21.175 ;
        RECT 77.085 17.010 81.895 17.085 ;
        RECT 82.215 17.010 82.710 21.855 ;
        RECT 84.240 21.855 90.680 22.350 ;
        RECT 84.240 17.010 84.735 21.855 ;
        RECT 85.055 21.175 89.865 21.535 ;
        RECT 85.055 17.085 85.415 21.175 ;
        RECT 85.725 17.395 89.195 20.865 ;
        RECT 89.505 17.085 89.865 21.175 ;
        RECT 85.055 17.010 89.865 17.085 ;
        RECT 90.185 17.010 90.680 21.855 ;
        RECT 95.710 17.830 96.670 27.120 ;
        RECT 97.630 25.520 99.230 25.920 ;
        RECT 96.990 24.320 97.310 25.520 ;
        RECT 98.270 24.720 99.870 25.120 ;
        RECT 100.190 24.320 100.510 25.520 ;
        RECT 97.630 23.920 99.230 24.320 ;
        RECT 97.750 18.560 98.590 22.180 ;
        RECT 100.830 18.560 101.790 27.120 ;
        RECT 103.150 18.560 104.470 20.690 ;
        RECT 105.580 18.560 107.570 34.390 ;
        RECT 108.690 32.430 110.130 33.630 ;
        RECT 109.770 28.830 110.130 32.430 ;
        RECT 110.850 32.430 112.290 33.630 ;
        RECT 110.850 28.830 111.210 32.430 ;
        RECT 111.930 28.830 112.290 32.430 ;
        RECT 113.010 32.430 114.450 33.630 ;
        RECT 113.010 28.830 113.370 32.430 ;
        RECT 114.090 28.830 114.450 32.430 ;
        RECT 115.170 32.430 116.610 33.630 ;
        RECT 115.170 28.830 115.530 32.430 ;
        RECT 116.250 28.830 116.610 32.430 ;
        RECT 117.330 32.430 118.770 33.630 ;
        RECT 117.330 28.830 117.690 32.430 ;
        RECT 118.410 28.830 118.770 32.430 ;
        RECT 119.490 32.430 120.930 33.630 ;
        RECT 119.490 28.830 119.850 32.430 ;
        RECT 120.570 28.830 120.930 32.430 ;
        RECT 121.650 32.430 123.090 33.630 ;
        RECT 121.650 28.830 122.010 32.430 ;
        RECT 122.730 28.830 123.090 32.430 ;
        RECT 123.810 32.430 125.250 33.630 ;
        RECT 123.810 28.830 124.170 32.430 ;
        RECT 124.890 28.830 125.250 32.430 ;
        RECT 125.970 32.430 127.410 33.630 ;
        RECT 125.970 28.830 126.330 32.430 ;
        RECT 109.770 19.230 111.210 21.630 ;
        RECT 111.930 19.230 113.370 21.630 ;
        RECT 114.090 19.230 115.530 21.630 ;
        RECT 116.250 19.230 117.690 21.630 ;
        RECT 118.410 19.230 119.850 21.630 ;
        RECT 120.570 19.230 122.010 21.630 ;
        RECT 122.730 19.230 124.170 21.630 ;
        RECT 124.890 19.230 126.330 21.630 ;
        RECT 128.590 18.560 129.150 34.390 ;
        RECT 131.480 26.770 132.440 33.760 ;
        RECT 133.400 32.960 135.640 33.360 ;
        RECT 132.760 30.960 133.080 32.160 ;
        RECT 134.040 31.360 136.280 31.760 ;
        RECT 136.600 30.960 136.920 32.160 ;
        RECT 133.400 29.760 135.640 30.160 ;
        RECT 133.400 26.770 134.360 28.650 ;
        RECT 137.240 26.770 138.200 33.760 ;
        RECT 141.400 26.770 142.360 33.750 ;
        RECT 143.320 32.950 145.560 33.350 ;
        RECT 142.680 30.950 143.000 32.150 ;
        RECT 143.960 31.350 146.200 31.750 ;
        RECT 146.520 30.950 146.840 32.150 ;
        RECT 143.320 29.750 145.560 30.150 ;
        RECT 143.320 26.770 144.280 28.770 ;
        RECT 147.160 26.770 148.120 33.750 ;
        RECT 131.480 26.760 148.120 26.770 ;
        RECT 131.320 26.740 148.120 26.760 ;
        RECT 150.840 26.740 159.410 76.910 ;
        RECT 131.320 20.020 159.410 26.740 ;
        RECT 131.320 18.560 159.390 20.020 ;
        RECT 0.580 15.920 90.680 17.010 ;
        RECT 0.580 8.910 64.420 15.920 ;
        RECT 68.300 15.910 74.740 15.920 ;
        RECT 76.270 15.910 82.710 15.920 ;
        RECT 84.240 15.910 90.680 15.920 ;
        RECT 68.300 13.755 74.740 14.250 ;
        RECT 68.300 8.910 68.795 13.755 ;
        RECT 69.115 13.075 73.925 13.435 ;
        RECT 69.115 8.985 69.475 13.075 ;
        RECT 69.785 9.295 73.255 12.765 ;
        RECT 73.565 8.985 73.925 13.075 ;
        RECT 69.115 8.910 73.925 8.985 ;
        RECT 74.245 8.910 74.740 13.755 ;
        RECT 76.270 13.755 82.710 14.250 ;
        RECT 76.270 8.910 76.765 13.755 ;
        RECT 77.085 13.075 81.895 13.435 ;
        RECT 77.085 8.985 77.445 13.075 ;
        RECT 77.755 9.295 81.225 12.765 ;
        RECT 81.535 8.985 81.895 13.075 ;
        RECT 77.085 8.910 81.895 8.985 ;
        RECT 82.215 8.910 82.710 13.755 ;
        RECT 84.240 13.755 90.680 14.250 ;
        RECT 84.240 8.910 84.735 13.755 ;
        RECT 85.055 13.075 89.865 13.435 ;
        RECT 85.055 8.985 85.415 13.075 ;
        RECT 85.725 9.295 89.195 12.765 ;
        RECT 89.505 8.985 89.865 13.075 ;
        RECT 85.055 8.910 89.865 8.985 ;
        RECT 90.185 8.910 90.680 13.755 ;
        RECT 0.580 8.860 90.680 8.910 ;
        RECT 97.120 8.860 159.390 18.560 ;
        RECT 0.580 7.760 159.390 8.860 ;
        RECT 0.580 7.600 153.290 7.760 ;
        RECT 0.610 7.320 153.290 7.600 ;
        RECT 0.610 7.250 4.640 7.320 ;
        RECT 64.030 7.230 98.700 7.320 ;
      LAYER met1 ;
        RECT 12.890 157.210 13.190 217.820 ;
        RECT 14.240 160.790 14.540 219.410 ;
        RECT 15.850 218.460 16.210 218.760 ;
        RECT 14.180 160.320 14.720 160.790 ;
        RECT 12.890 156.850 13.210 157.210 ;
        RECT 12.890 156.760 13.190 156.850 ;
        RECT 15.880 152.450 16.180 218.460 ;
        RECT 19.570 164.980 19.870 220.990 ;
        RECT 20.390 168.250 20.690 220.130 ;
        RECT 21.080 167.570 21.380 223.550 ;
        RECT 56.765 213.100 58.570 213.130 ;
        RECT 56.765 212.290 60.880 213.100 ;
        RECT 54.000 211.890 150.000 212.290 ;
        RECT 54.000 211.770 150.100 211.890 ;
        RECT 53.860 210.290 150.100 211.770 ;
        RECT 53.220 189.770 53.540 209.230 ;
        RECT 53.860 191.130 54.820 210.290 ;
        RECT 55.780 189.770 56.740 209.230 ;
        RECT 62.220 189.770 62.540 208.730 ;
        RECT 62.860 191.130 63.820 210.290 ;
        RECT 64.780 205.780 65.740 208.730 ;
        RECT 64.770 193.760 65.750 205.780 ;
        RECT 64.780 189.770 65.740 193.760 ;
        RECT 71.220 189.770 71.540 208.730 ;
        RECT 71.860 191.130 72.820 210.290 ;
        RECT 73.780 189.770 74.740 208.730 ;
        RECT 80.220 189.770 80.540 208.730 ;
        RECT 80.860 191.130 81.820 210.290 ;
        RECT 82.780 189.770 83.740 208.730 ;
        RECT 89.220 201.610 89.540 201.730 ;
        RECT 88.900 189.770 89.540 201.610 ;
        RECT 89.860 198.130 90.820 210.290 ;
        RECT 53.020 189.130 89.540 189.770 ;
        RECT 53.020 188.810 89.480 189.130 ;
        RECT 73.840 187.190 75.040 188.810 ;
        RECT 91.780 187.830 92.740 201.730 ;
        RECT 98.220 188.950 98.540 208.730 ;
        RECT 98.860 191.130 99.820 210.290 ;
        RECT 100.780 204.270 101.740 208.730 ;
        RECT 100.750 203.310 101.770 204.270 ;
        RECT 100.780 195.780 101.740 201.730 ;
        RECT 91.050 187.770 92.740 187.830 ;
        RECT 95.340 188.630 98.540 188.950 ;
        RECT 100.780 188.780 101.740 194.730 ;
        RECT 54.900 185.790 57.600 187.190 ;
        RECT 73.700 185.790 75.200 187.190 ;
        RECT 80.860 186.810 92.780 187.770 ;
        RECT 20.110 167.270 21.380 167.570 ;
        RECT 19.540 164.680 19.900 164.980 ;
        RECT 20.110 164.120 20.410 167.270 ;
        RECT 20.590 165.680 21.470 166.020 ;
        RECT 20.060 163.790 20.410 164.120 ;
        RECT 21.820 164.070 22.120 168.610 ;
        RECT 22.690 167.350 22.990 170.060 ;
        RECT 23.290 165.680 24.170 166.020 ;
        RECT 20.060 162.010 20.360 163.790 ;
        RECT 20.590 163.280 21.470 163.620 ;
        RECT 23.290 163.280 24.170 163.620 ;
        RECT 26.300 162.580 26.620 163.030 ;
        RECT 25.520 162.260 26.620 162.580 ;
        RECT 20.000 161.710 20.420 162.010 ;
        RECT 20.590 160.880 21.470 161.220 ;
        RECT 23.290 160.880 24.170 161.220 ;
        RECT 18.790 160.700 19.090 160.760 ;
        RECT 18.400 160.400 19.090 160.700 ;
        RECT 18.790 160.340 19.090 160.400 ;
        RECT 20.590 159.280 21.470 159.620 ;
        RECT 23.290 159.280 24.170 159.620 ;
        RECT 20.590 157.680 21.470 158.020 ;
        RECT 25.295 157.970 26.480 158.305 ;
        RECT 26.145 157.530 26.480 157.970 ;
        RECT 19.940 157.180 20.240 157.240 ;
        RECT 26.115 157.195 26.510 157.530 ;
        RECT 19.190 156.880 20.240 157.180 ;
        RECT 19.940 156.820 20.240 156.880 ;
        RECT 20.590 156.080 21.470 156.420 ;
        RECT 23.290 156.080 24.170 156.420 ;
        RECT 20.590 154.480 21.470 154.820 ;
        RECT 23.290 154.480 24.170 154.820 ;
        RECT 25.600 154.390 25.900 154.450 ;
        RECT 25.600 154.090 26.360 154.390 ;
        RECT 25.600 154.030 25.900 154.090 ;
        RECT 20.590 152.880 21.470 153.220 ;
        RECT 23.290 152.880 24.170 153.220 ;
        RECT 18.860 152.780 19.160 152.840 ;
        RECT 18.280 152.480 19.160 152.780 ;
        RECT 18.860 152.420 19.160 152.480 ;
        RECT 20.590 151.280 21.470 151.620 ;
        RECT 23.290 151.280 24.170 151.620 ;
        RECT 20.590 150.480 21.470 150.820 ;
        RECT 23.290 150.480 24.170 150.820 ;
        RECT 6.160 139.980 8.160 140.010 ;
        RECT 6.160 137.980 11.830 139.980 ;
        RECT 20.560 138.530 23.040 139.410 ;
        RECT 6.160 137.950 8.160 137.980 ;
        RECT 28.780 109.720 30.000 160.920 ;
        RECT 32.690 157.840 33.650 158.850 ;
        RECT 32.660 156.880 33.680 157.840 ;
        RECT 32.690 111.890 33.650 156.880 ;
        RECT 49.250 135.950 49.570 163.030 ;
        RECT 50.260 135.560 50.560 170.060 ;
        RECT 54.900 169.190 56.100 185.790 ;
        RECT 80.220 175.130 80.540 186.480 ;
        RECT 80.860 175.130 81.820 186.810 ;
        RECT 82.780 173.770 83.740 186.230 ;
        RECT 89.220 175.130 89.540 186.480 ;
        RECT 89.860 175.130 90.820 186.810 ;
        RECT 91.050 186.750 92.010 186.810 ;
        RECT 80.020 172.810 89.980 173.770 ;
        RECT 91.780 173.450 92.740 185.730 ;
        RECT 95.340 173.450 95.660 188.630 ;
        RECT 91.780 172.930 95.660 173.450 ;
        RECT 54.900 167.790 57.600 169.190 ;
        RECT 80.220 162.130 80.540 172.810 ;
        RECT 80.860 161.760 81.820 170.730 ;
        RECT 82.780 162.130 83.740 172.810 ;
        RECT 89.220 162.130 89.540 172.810 ;
        RECT 85.990 161.770 86.950 161.830 ;
        RECT 89.860 161.770 90.820 170.730 ;
        RECT 91.780 162.130 92.740 172.930 ;
        RECT 95.340 166.450 95.660 172.930 ;
        RECT 95.340 166.130 97.690 166.450 ;
        RECT 85.080 161.760 90.820 161.770 ;
        RECT 80.860 160.820 90.820 161.760 ;
        RECT 80.860 160.810 81.820 160.820 ;
        RECT 85.080 160.810 90.820 160.820 ;
        RECT 85.990 160.750 86.950 160.810 ;
        RECT 77.370 158.950 78.630 160.150 ;
        RECT 103.000 159.570 105.000 210.290 ;
        RECT 108.260 187.830 109.220 201.730 ;
        RECT 110.180 198.130 111.140 210.290 ;
        RECT 111.460 201.610 111.780 201.730 ;
        RECT 111.460 189.770 112.100 201.610 ;
        RECT 117.260 189.770 118.220 208.730 ;
        RECT 119.180 191.130 120.140 210.290 ;
        RECT 120.460 189.770 120.780 208.730 ;
        RECT 126.260 189.770 127.220 208.730 ;
        RECT 128.180 191.130 129.140 210.290 ;
        RECT 129.460 189.770 129.780 208.730 ;
        RECT 135.260 205.780 136.220 208.730 ;
        RECT 135.250 193.760 136.230 205.780 ;
        RECT 135.260 189.770 136.220 193.760 ;
        RECT 137.180 191.130 138.140 210.290 ;
        RECT 138.460 189.770 138.780 208.730 ;
        RECT 144.260 189.770 145.220 209.230 ;
        RECT 146.180 191.130 147.140 210.290 ;
        RECT 148.900 210.090 150.100 210.290 ;
        RECT 152.200 210.090 153.600 210.190 ;
        RECT 147.460 189.770 147.780 209.230 ;
        RECT 148.900 208.890 153.600 210.090 ;
        RECT 152.200 208.790 153.600 208.890 ;
        RECT 156.800 208.790 159.100 210.190 ;
        RECT 157.900 192.190 159.100 208.790 ;
        RECT 151.400 190.790 153.600 192.190 ;
        RECT 156.800 190.790 159.100 192.190 ;
        RECT 111.460 189.130 147.980 189.770 ;
        RECT 111.520 188.810 147.980 189.130 ;
        RECT 108.260 187.770 109.950 187.830 ;
        RECT 108.220 186.810 120.140 187.770 ;
        RECT 125.960 187.190 127.160 188.810 ;
        RECT 108.990 186.750 109.950 186.810 ;
        RECT 108.260 173.340 109.220 185.730 ;
        RECT 110.180 175.130 111.140 186.810 ;
        RECT 111.460 175.130 111.780 186.480 ;
        RECT 117.260 173.770 118.220 186.230 ;
        RECT 119.180 175.130 120.140 186.810 ;
        RECT 120.460 175.130 120.780 186.480 ;
        RECT 125.800 185.790 127.300 187.190 ;
        RECT 143.400 185.790 146.100 187.190 ;
        RECT 105.750 173.040 109.220 173.340 ;
        RECT 105.750 160.240 106.050 173.040 ;
        RECT 108.260 162.130 109.220 173.040 ;
        RECT 111.020 172.810 120.980 173.770 ;
        RECT 110.180 161.770 111.140 170.730 ;
        RECT 111.460 162.130 111.780 172.810 ;
        RECT 117.260 162.130 118.220 172.810 ;
        RECT 114.050 161.770 115.010 161.830 ;
        RECT 110.180 161.760 115.920 161.770 ;
        RECT 119.180 161.760 120.140 170.730 ;
        RECT 120.460 162.130 120.780 172.810 ;
        RECT 144.900 169.190 146.100 185.790 ;
        RECT 151.400 174.150 152.600 190.790 ;
        RECT 158.080 174.150 159.100 176.130 ;
        RECT 151.400 172.890 153.490 174.150 ;
        RECT 152.290 172.830 153.490 172.890 ;
        RECT 156.910 172.830 159.100 174.150 ;
        RECT 143.400 167.790 146.100 169.190 ;
        RECT 110.180 160.820 120.140 161.760 ;
        RECT 110.180 160.810 115.920 160.820 ;
        RECT 119.180 160.810 120.140 160.820 ;
        RECT 114.050 160.750 115.010 160.810 ;
        RECT 105.750 159.940 114.080 160.240 ;
        RECT 55.400 149.790 57.600 151.190 ;
        RECT 73.870 151.090 75.070 151.150 ;
        RECT 77.400 151.090 78.600 158.950 ;
        RECT 103.000 158.610 107.310 159.570 ;
        RECT 92.650 158.340 92.950 158.370 ;
        RECT 91.420 158.040 92.950 158.340 ;
        RECT 92.650 158.010 92.950 158.040 ;
        RECT 73.870 149.890 78.600 151.090 ;
        RECT 81.100 152.990 100.600 156.390 ;
        RECT 103.000 156.290 105.000 158.610 ;
        RECT 107.420 155.910 107.720 158.500 ;
        RECT 108.220 157.340 109.100 157.680 ;
        RECT 110.920 157.340 111.800 157.680 ;
        RECT 113.780 156.880 114.080 159.940 ;
        RECT 112.560 156.230 113.440 156.260 ;
        RECT 112.560 155.350 116.670 156.230 ;
        RECT 157.900 156.150 159.100 172.830 ;
        RECT 112.560 155.320 113.440 155.350 ;
        RECT 156.910 154.890 159.100 156.150 ;
        RECT 156.910 154.830 158.110 154.890 ;
        RECT 109.320 153.940 109.620 154.000 ;
        RECT 106.820 153.640 109.620 153.940 ;
        RECT 109.320 153.580 109.620 153.640 ;
        RECT 110.100 153.340 110.980 153.380 ;
        RECT 110.100 153.040 111.600 153.340 ;
        RECT 73.870 149.830 75.070 149.890 ;
        RECT 50.230 135.260 50.590 135.560 ;
        RECT 55.400 133.190 56.600 149.790 ;
        RECT 81.100 140.290 84.500 152.990 ;
        RECT 90.400 148.165 91.600 150.920 ;
        RECT 89.325 145.115 92.375 148.165 ;
        RECT 97.300 140.290 100.600 152.990 ;
        RECT 107.400 152.240 108.280 152.580 ;
        RECT 110.100 152.240 110.980 152.580 ;
        RECT 107.400 151.740 108.280 151.780 ;
        RECT 107.400 151.440 108.900 151.740 ;
        RECT 105.600 151.040 106.480 151.380 ;
        RECT 105.600 149.740 106.480 149.780 ;
        RECT 81.100 136.990 100.600 140.290 ;
        RECT 105.000 149.440 106.480 149.740 ;
        RECT 105.000 137.740 105.300 149.440 ;
        RECT 107.400 149.040 108.280 149.380 ;
        RECT 107.400 148.540 108.280 148.580 ;
        RECT 108.600 148.540 108.900 151.440 ;
        RECT 111.300 150.540 111.600 153.040 ;
        RECT 144.370 152.390 145.570 152.450 ;
        RECT 142.370 151.190 145.570 152.390 ;
        RECT 144.370 151.130 145.570 151.190 ;
        RECT 111.900 150.540 112.780 150.580 ;
        RECT 111.300 150.240 112.780 150.540 ;
        RECT 110.100 149.840 110.980 150.180 ;
        RECT 107.400 148.240 108.900 148.540 ;
        RECT 111.900 148.140 112.780 148.180 ;
        RECT 111.900 147.840 113.400 148.140 ;
        RECT 111.900 147.340 112.780 147.380 ;
        RECT 111.300 147.040 112.780 147.340 ;
        RECT 107.400 146.640 108.280 146.980 ;
        RECT 110.100 146.640 110.980 146.980 ;
        RECT 110.100 146.140 110.980 146.180 ;
        RECT 111.300 146.140 111.600 147.040 ;
        RECT 110.100 145.840 111.600 146.140 ;
        RECT 105.600 145.740 106.480 145.780 ;
        RECT 105.600 145.440 107.100 145.740 ;
        RECT 106.800 144.540 107.100 145.440 ;
        RECT 107.400 145.040 108.280 145.380 ;
        RECT 110.100 145.040 110.980 145.380 ;
        RECT 107.400 144.540 108.280 144.580 ;
        RECT 106.800 144.240 108.280 144.540 ;
        RECT 111.300 143.340 111.600 145.840 ;
        RECT 111.900 144.140 112.780 144.180 ;
        RECT 113.100 144.140 113.400 147.840 ;
        RECT 111.900 143.840 113.400 144.140 ;
        RECT 111.900 143.340 112.780 143.380 ;
        RECT 111.300 143.040 112.780 143.340 ;
        RECT 107.400 142.640 108.280 142.980 ;
        RECT 110.100 142.640 110.980 142.980 ;
        RECT 105.600 141.740 106.480 141.780 ;
        RECT 105.600 141.440 106.500 141.740 ;
        RECT 106.200 141.140 107.100 141.440 ;
        RECT 106.800 138.140 107.100 141.140 ;
        RECT 107.400 140.240 108.280 140.580 ;
        RECT 110.100 140.240 110.980 140.580 ;
        RECT 112.290 140.110 112.710 140.410 ;
        RECT 112.350 139.610 112.650 140.110 ;
        RECT 107.400 138.640 108.280 138.980 ;
        RECT 110.100 138.640 110.980 138.980 ;
        RECT 107.400 138.140 108.280 138.180 ;
        RECT 106.800 137.840 108.280 138.140 ;
        RECT 110.100 137.840 110.980 138.180 ;
        RECT 105.600 137.740 106.480 137.780 ;
        RECT 105.000 137.440 106.480 137.740 ;
        RECT 97.840 133.190 99.040 136.990 ;
        RECT 105.000 134.040 105.300 137.440 ;
        RECT 110.100 137.340 110.980 137.380 ;
        RECT 113.100 137.340 113.400 143.840 ;
        RECT 110.100 137.040 113.400 137.340 ;
        RECT 107.400 136.240 108.280 136.580 ;
        RECT 110.100 136.240 110.980 136.580 ;
        RECT 105.730 135.910 106.150 136.210 ;
        RECT 105.790 135.370 106.090 135.910 ;
        RECT 107.400 135.440 108.280 135.780 ;
        RECT 110.100 135.440 110.980 135.780 ;
        RECT 107.400 134.640 108.280 134.980 ;
        RECT 110.100 134.640 110.980 134.980 ;
        RECT 105.000 133.740 111.480 134.040 ;
        RECT 55.400 131.790 57.700 133.190 ;
        RECT 73.800 133.090 75.100 133.190 ;
        RECT 80.200 133.090 81.600 133.190 ;
        RECT 73.800 131.890 81.600 133.090 ;
        RECT 73.800 131.790 75.100 131.890 ;
        RECT 80.200 131.790 81.600 131.890 ;
        RECT 97.800 131.790 99.100 133.190 ;
        RECT 102.650 132.640 103.100 133.090 ;
        RECT 102.720 124.630 103.040 132.640 ;
        RECT 103.360 123.280 104.320 133.030 ;
        RECT 104.640 132.070 108.910 133.030 ;
        RECT 104.640 124.630 105.600 132.070 ;
        RECT 108.180 129.040 109.120 129.920 ;
        RECT 108.210 127.510 109.090 129.040 ;
        RECT 25.580 103.150 154.620 108.400 ;
        RECT 25.580 75.310 53.920 103.150 ;
        RECT 74.290 102.400 75.250 103.150 ;
        RECT 74.230 101.440 75.310 102.400 ;
        RECT 75.570 98.880 75.890 100.700 ;
        RECT 75.570 97.100 75.900 98.880 ;
        RECT 75.580 96.540 75.900 97.100 ;
        RECT 76.210 96.540 77.170 103.150 ;
        RECT 80.050 102.400 81.010 103.150 ;
        RECT 79.990 101.440 81.070 102.400 ;
        RECT 83.650 101.000 89.890 103.150 ;
        RECT 113.030 101.160 114.230 101.220 ;
        RECT 109.080 101.140 114.230 101.160 ;
        RECT 102.410 101.080 103.610 101.140 ;
        RECT 91.760 101.000 92.960 101.060 ;
        RECT 78.130 99.750 79.090 100.700 ;
        RECT 83.630 99.800 92.960 101.000 ;
        RECT 78.130 97.100 79.100 99.750 ;
        RECT 78.140 96.540 79.100 97.100 ;
        RECT 64.410 90.650 64.730 94.780 ;
        RECT 65.050 94.700 66.010 94.780 ;
        RECT 65.050 91.180 66.040 94.700 ;
        RECT 66.970 93.880 67.930 94.780 ;
        RECT 66.970 91.180 67.960 93.880 ;
        RECT 75.550 92.940 75.900 96.540 ;
        RECT 76.190 92.940 77.170 96.540 ;
        RECT 78.110 92.940 79.100 96.540 ;
        RECT 65.080 90.650 66.040 91.180 ;
        RECT 67.000 90.650 67.960 91.180 ;
        RECT 64.400 87.050 64.730 90.650 ;
        RECT 65.040 87.050 66.040 90.650 ;
        RECT 66.960 87.050 67.960 90.650 ;
        RECT 75.580 92.550 75.900 92.940 ;
        RECT 76.210 92.550 77.170 92.940 ;
        RECT 78.140 92.550 79.100 92.940 ;
        RECT 75.580 88.950 75.910 92.550 ;
        RECT 76.210 88.950 77.190 92.550 ;
        RECT 78.140 88.950 79.110 92.550 ;
        RECT 75.580 88.390 75.900 88.950 ;
        RECT 76.210 88.390 77.170 88.950 ;
        RECT 78.140 88.390 79.100 88.950 ;
        RECT 64.410 86.650 64.730 87.050 ;
        RECT 65.080 86.650 66.040 87.050 ;
        RECT 67.000 86.650 67.960 87.050 ;
        RECT 64.410 83.050 64.750 86.650 ;
        RECT 65.070 83.050 66.040 86.650 ;
        RECT 66.990 83.050 67.960 86.650 ;
        RECT 75.550 84.790 75.900 88.390 ;
        RECT 76.190 84.790 77.170 88.390 ;
        RECT 78.110 84.790 79.100 88.390 ;
        RECT 75.580 84.390 75.900 84.790 ;
        RECT 64.410 82.520 64.730 83.050 ;
        RECT 65.080 82.520 66.040 83.050 ;
        RECT 67.000 82.520 67.960 83.050 ;
        RECT 64.410 78.920 64.740 82.520 ;
        RECT 65.060 78.920 66.040 82.520 ;
        RECT 66.980 78.920 67.960 82.520 ;
        RECT 75.570 80.790 75.900 84.390 ;
        RECT 75.580 80.230 75.900 80.790 ;
        RECT 76.210 80.230 77.170 84.790 ;
        RECT 78.140 84.390 79.100 84.790 ;
        RECT 78.130 80.790 79.100 84.390 ;
        RECT 78.140 80.230 79.100 80.790 ;
        RECT 64.410 78.530 64.730 78.920 ;
        RECT 65.080 78.530 66.040 78.920 ;
        RECT 67.000 78.530 67.960 78.920 ;
        RECT 39.680 73.700 53.880 75.310 ;
        RECT 39.400 72.580 53.880 73.700 ;
        RECT 39.400 72.520 40.460 72.580 ;
        RECT 24.050 72.230 25.250 72.290 ;
        RECT 37.730 72.230 38.690 72.240 ;
        RECT 6.440 71.000 7.760 72.200 ;
        RECT 24.050 71.030 38.690 72.230 ;
        RECT 6.500 59.560 7.700 71.000 ;
        RECT 24.050 70.970 25.250 71.030 ;
        RECT 35.170 69.140 35.490 71.030 ;
        RECT 35.810 69.140 36.770 70.670 ;
        RECT 37.730 69.140 38.690 71.030 ;
        RECT 35.160 68.400 35.490 69.140 ;
        RECT 35.160 66.010 35.480 68.400 ;
        RECT 35.800 67.470 36.770 69.140 ;
        RECT 37.720 67.830 38.690 69.140 ;
        RECT 35.800 66.460 36.760 67.470 ;
        RECT 35.160 65.540 35.510 66.010 ;
        RECT 35.800 65.540 36.790 66.460 ;
        RECT 37.720 65.540 38.680 67.830 ;
        RECT 35.190 64.120 35.510 65.540 ;
        RECT 35.830 64.120 36.790 65.540 ;
        RECT 46.550 64.650 53.880 72.580 ;
        RECT 64.410 74.930 64.750 78.530 ;
        RECT 65.070 74.930 66.040 78.530 ;
        RECT 66.990 74.930 67.960 78.530 ;
        RECT 75.550 76.630 75.900 80.230 ;
        RECT 76.190 76.630 77.170 80.230 ;
        RECT 78.110 76.630 79.100 80.230 ;
        RECT 75.580 76.100 75.900 76.630 ;
        RECT 64.410 74.400 64.730 74.930 ;
        RECT 65.080 74.400 66.040 74.930 ;
        RECT 67.000 74.400 67.960 74.930 ;
        RECT 64.410 70.800 64.740 74.400 ;
        RECT 65.060 70.800 66.040 74.400 ;
        RECT 66.980 70.800 67.960 74.400 ;
        RECT 75.570 72.500 75.900 76.100 ;
        RECT 64.410 70.390 64.730 70.800 ;
        RECT 65.080 70.390 66.040 70.800 ;
        RECT 67.000 70.390 67.960 70.800 ;
        RECT 64.410 66.790 64.770 70.390 ;
        RECT 65.080 66.790 66.050 70.390 ;
        RECT 67.000 66.790 67.970 70.390 ;
        RECT 75.580 67.810 75.900 72.500 ;
        RECT 76.210 71.940 77.170 76.630 ;
        RECT 78.140 76.100 79.100 76.630 ;
        RECT 78.130 72.500 79.100 76.100 ;
        RECT 76.210 68.340 77.180 71.940 ;
        RECT 76.210 67.810 77.170 68.340 ;
        RECT 78.140 67.810 79.100 72.500 ;
        RECT 64.410 66.260 64.730 66.790 ;
        RECT 35.180 62.890 35.510 64.120 ;
        RECT 35.180 60.520 35.500 62.890 ;
        RECT 35.820 62.010 36.790 64.120 ;
        RECT 35.820 60.520 36.780 62.010 ;
        RECT 37.740 60.980 38.700 64.120 ;
        RECT 46.480 61.120 61.210 64.650 ;
        RECT 64.410 62.660 64.760 66.260 ;
        RECT 64.410 62.270 64.730 62.660 ;
        RECT 65.080 62.270 66.040 66.790 ;
        RECT 67.000 62.270 67.960 66.790 ;
        RECT 75.560 64.210 75.900 67.810 ;
        RECT 76.200 64.210 77.170 67.810 ;
        RECT 78.120 64.210 79.100 67.810 ;
        RECT 83.650 67.100 89.890 99.800 ;
        RECT 91.760 99.740 92.960 99.800 ;
        RECT 97.530 101.000 98.730 101.060 ;
        RECT 99.430 101.000 103.610 101.080 ;
        RECT 97.530 99.880 103.610 101.000 ;
        RECT 97.530 99.800 101.390 99.880 ;
        RECT 102.410 99.820 103.610 99.880 ;
        RECT 108.310 99.960 114.230 101.140 ;
        RECT 108.310 99.880 112.370 99.960 ;
        RECT 113.030 99.900 114.230 99.960 ;
        RECT 118.930 101.160 120.130 101.220 ;
        RECT 118.930 99.960 122.930 101.160 ;
        RECT 118.930 99.900 120.130 99.960 ;
        RECT 108.310 99.820 109.510 99.880 ;
        RECT 97.530 99.740 98.730 99.800 ;
        RECT 111.115 82.075 111.445 99.880 ;
        RECT 121.730 85.120 122.930 99.960 ;
        RECT 121.700 83.920 122.960 85.120 ;
        RECT 111.085 81.745 111.475 82.075 ;
        RECT 135.180 73.460 139.660 103.150 ;
        RECT 158.460 96.210 159.420 112.910 ;
        RECT 150.810 95.250 159.420 96.210 ;
        RECT 138.520 73.430 139.580 73.460 ;
        RECT 126.400 68.690 127.600 68.750 ;
        RECT 140.080 68.690 141.040 68.700 ;
        RECT 108.790 67.460 110.110 68.660 ;
        RECT 126.400 67.490 141.040 68.690 ;
        RECT 83.620 66.140 90.370 67.100 ;
        RECT 83.620 65.820 84.610 66.140 ;
        RECT 83.590 64.860 84.670 65.820 ;
        RECT 37.740 60.520 38.710 60.980 ;
        RECT 6.500 58.360 25.060 59.560 ;
        RECT 6.370 47.360 7.570 54.700 ;
        RECT 23.860 53.410 25.060 58.360 ;
        RECT 29.070 58.920 32.580 58.970 ;
        RECT 37.750 58.920 38.710 60.520 ;
        RECT 46.480 60.060 61.350 61.120 ;
        RECT 44.770 58.940 45.730 59.000 ;
        RECT 40.250 58.920 45.730 58.940 ;
        RECT 29.070 58.010 45.730 58.920 ;
        RECT 31.050 57.980 45.730 58.010 ;
        RECT 31.050 57.960 41.950 57.980 ;
        RECT 27.755 48.770 28.085 48.800 ;
        RECT 30.410 48.770 30.730 57.070 ;
        RECT 31.050 48.770 32.010 57.960 ;
        RECT 34.830 57.940 35.910 57.960 ;
        RECT 38.980 57.940 40.060 57.960 ;
        RECT 40.990 57.110 41.950 57.960 ;
        RECT 44.770 57.920 45.730 57.980 ;
        RECT 32.970 54.800 33.930 57.070 ;
        RECT 27.705 48.440 30.730 48.770 ;
        RECT 27.755 48.410 28.085 48.440 ;
        RECT 6.370 46.160 25.020 47.360 ;
        RECT 6.280 35.940 7.600 37.140 ;
        RECT 23.820 35.950 25.020 46.160 ;
        RECT 30.400 45.170 30.730 48.440 ;
        RECT 31.040 45.170 32.010 48.770 ;
        RECT 30.410 44.660 30.730 45.170 ;
        RECT 31.050 44.660 32.010 45.170 ;
        RECT 30.400 44.060 30.730 44.660 ;
        RECT 30.400 41.060 30.720 44.060 ;
        RECT 31.040 42.790 32.010 44.660 ;
        RECT 32.960 53.470 33.930 54.800 ;
        RECT 32.960 52.960 33.920 53.470 ;
        RECT 32.960 49.360 33.930 52.960 ;
        RECT 37.755 49.485 38.145 49.815 ;
        RECT 31.040 41.060 32.000 42.790 ;
        RECT 32.960 38.880 33.920 49.360 ;
        RECT 37.785 48.810 38.115 49.485 ;
        RECT 40.320 48.810 40.640 57.110 ;
        RECT 40.960 55.770 41.950 57.110 ;
        RECT 40.960 54.570 41.920 55.770 ;
        RECT 37.615 48.480 40.640 48.810 ;
        RECT 40.310 45.210 40.640 48.480 ;
        RECT 40.320 44.700 40.640 45.210 ;
        RECT 40.310 44.230 40.640 44.700 ;
        RECT 40.950 53.510 41.920 54.570 ;
        RECT 40.950 53.000 41.910 53.510 ;
        RECT 40.950 49.400 41.920 53.000 ;
        RECT 40.310 41.100 40.630 44.230 ;
        RECT 40.950 41.100 41.910 49.400 ;
        RECT 42.880 48.810 43.840 57.110 ;
        RECT 42.870 45.210 43.840 48.810 ;
        RECT 46.550 45.990 53.880 60.060 ;
        RECT 55.940 53.660 56.260 58.830 ;
        RECT 56.580 55.230 57.540 60.060 ;
        RECT 60.390 60.040 61.350 60.060 ;
        RECT 58.500 52.180 59.460 58.830 ;
        RECT 64.410 58.670 64.770 62.270 ;
        RECT 65.080 58.670 66.050 62.270 ;
        RECT 67.000 58.670 67.970 62.270 ;
        RECT 75.580 59.230 75.900 64.210 ;
        RECT 76.210 63.650 77.170 64.210 ;
        RECT 76.210 61.400 77.180 63.650 ;
        RECT 76.220 60.050 77.180 61.400 ;
        RECT 78.140 59.430 79.100 64.210 ;
        RECT 84.930 59.430 85.250 63.650 ;
        RECT 85.570 60.050 86.530 66.140 ;
        RECT 89.410 65.790 90.370 66.140 ;
        RECT 89.350 64.830 90.430 65.790 ;
        RECT 78.140 59.230 85.250 59.430 ;
        RECT 75.580 58.910 85.250 59.230 ;
        RECT 64.410 58.140 64.730 58.670 ;
        RECT 64.410 55.000 64.760 58.140 ;
        RECT 64.440 52.180 64.760 55.000 ;
        RECT 65.080 53.380 66.040 58.670 ;
        RECT 65.050 52.420 66.070 53.380 ;
        RECT 67.000 52.290 67.960 58.670 ;
        RECT 78.140 58.470 85.250 58.910 ;
        RECT 78.140 58.130 79.100 58.470 ;
        RECT 75.510 52.290 75.830 58.130 ;
        RECT 76.150 52.990 77.110 58.130 ;
        RECT 78.070 56.120 79.100 58.130 ;
        RECT 87.490 56.295 88.450 63.650 ;
        RECT 104.235 56.295 104.565 56.325 ;
        RECT 78.070 54.530 79.030 56.120 ;
        RECT 87.425 55.965 104.565 56.295 ;
        RECT 87.490 55.390 88.450 55.965 ;
        RECT 104.235 55.935 104.565 55.965 ;
        RECT 108.850 56.020 110.050 67.460 ;
        RECT 126.400 67.430 127.600 67.490 ;
        RECT 137.520 65.600 137.840 67.490 ;
        RECT 138.160 65.600 139.120 67.130 ;
        RECT 140.080 65.600 141.040 67.490 ;
        RECT 137.510 64.860 137.840 65.600 ;
        RECT 137.510 62.470 137.830 64.860 ;
        RECT 138.150 63.930 139.120 65.600 ;
        RECT 140.070 64.290 141.040 65.600 ;
        RECT 138.150 62.920 139.110 63.930 ;
        RECT 137.510 62.000 137.860 62.470 ;
        RECT 138.150 62.000 139.140 62.920 ;
        RECT 140.070 62.000 141.030 64.290 ;
        RECT 137.540 60.580 137.860 62.000 ;
        RECT 138.180 60.580 139.140 62.000 ;
        RECT 137.530 59.350 137.860 60.580 ;
        RECT 137.530 56.980 137.850 59.350 ;
        RECT 138.170 58.470 139.140 60.580 ;
        RECT 138.170 56.980 139.130 58.470 ;
        RECT 140.090 57.440 141.050 60.580 ;
        RECT 140.090 56.980 141.060 57.440 ;
        RECT 108.850 54.820 127.410 56.020 ;
        RECT 88.090 53.750 92.540 54.100 ;
        RECT 88.090 53.430 97.310 53.750 ;
        RECT 88.090 52.880 92.540 53.430 ;
        RECT 67.000 52.180 75.950 52.290 ;
        RECT 58.500 51.330 75.950 52.180 ;
        RECT 58.500 51.250 67.960 51.330 ;
        RECT 58.540 51.220 67.960 51.250 ;
        RECT 71.900 49.890 73.100 49.950 ;
        RECT 64.170 49.225 73.100 49.890 ;
        RECT 63.010 48.895 73.100 49.225 ;
        RECT 64.150 48.690 73.100 48.895 ;
        RECT 60.310 45.990 61.270 46.000 ;
        RECT 46.550 45.440 63.200 45.990 ;
        RECT 42.880 44.700 43.840 45.210 ;
        RECT 46.670 45.030 63.200 45.440 ;
        RECT 42.870 43.170 43.840 44.700 ;
        RECT 52.580 43.550 53.540 45.030 ;
        RECT 60.310 44.790 61.270 45.030 ;
        RECT 62.230 44.990 63.200 45.030 ;
        RECT 60.250 43.830 61.330 44.790 ;
        RECT 42.870 39.230 43.830 43.170 ;
        RECT 61.590 40.080 61.910 43.220 ;
        RECT 62.230 41.370 63.190 44.990 ;
        RECT 61.590 39.620 61.920 40.080 ;
        RECT 62.230 39.620 63.200 41.370 ;
        RECT 64.150 39.620 65.110 48.690 ;
        RECT 71.900 48.630 73.100 48.690 ;
        RECT 77.830 49.890 79.030 49.950 ;
        RECT 77.830 49.880 80.670 49.890 ;
        RECT 81.620 49.880 82.820 49.940 ;
        RECT 77.830 48.680 82.820 49.880 ;
        RECT 77.830 48.630 79.030 48.680 ;
        RECT 81.620 48.620 82.820 48.680 ;
        RECT 30.410 38.830 34.000 38.880 ;
        RECT 30.410 38.560 40.650 38.830 ;
        RECT 6.340 20.170 7.540 35.940 ;
        RECT 30.410 33.300 30.730 38.560 ;
        RECT 32.960 38.510 40.650 38.560 ;
        RECT 32.960 36.900 33.920 38.510 ;
        RECT 31.050 31.200 32.010 36.900 ;
        RECT 32.960 34.900 33.930 36.900 ;
        RECT 32.970 33.300 33.930 34.900 ;
        RECT 40.330 33.290 40.650 38.510 ;
        RECT 42.870 38.270 57.320 39.230 ;
        RECT 42.870 36.890 43.830 38.270 ;
        RECT 40.970 31.320 41.930 36.890 ;
        RECT 42.870 35.020 43.850 36.890 ;
        RECT 42.890 33.290 43.850 35.020 ;
        RECT 57.000 35.190 57.320 38.270 ;
        RECT 61.600 35.190 61.920 39.620 ;
        RECT 62.240 35.500 63.200 39.620 ;
        RECT 57.000 34.870 61.920 35.190 ;
        RECT 61.600 33.340 61.920 34.870 ;
        RECT 64.160 24.190 65.120 39.100 ;
        RECT 69.995 27.920 73.045 28.755 ;
        RECT 77.965 27.920 81.015 28.755 ;
        RECT 85.935 27.920 88.985 28.755 ;
        RECT 91.790 27.920 92.990 49.870 ;
        RECT 69.995 26.720 92.990 27.920 ;
        RECT 69.995 25.705 73.045 26.720 ;
        RECT 77.965 25.705 81.015 26.720 ;
        RECT 85.935 25.705 88.985 26.720 ;
        RECT 64.160 23.230 79.870 24.190 ;
        RECT 78.910 20.655 79.870 23.230 ;
        RECT 4.630 19.620 5.190 19.680 ;
        RECT 6.340 19.620 30.200 20.170 ;
        RECT 4.630 19.060 30.200 19.620 ;
        RECT 4.630 19.000 5.190 19.060 ;
        RECT 6.340 18.970 30.200 19.060 ;
        RECT 69.995 17.605 73.045 20.655 ;
        RECT 77.965 17.605 81.015 20.655 ;
        RECT 85.935 20.370 88.985 20.655 ;
        RECT 91.790 20.370 92.990 26.720 ;
        RECT 96.990 23.120 97.310 53.430 ;
        RECT 108.720 43.820 109.920 51.160 ;
        RECT 126.210 49.870 127.410 54.820 ;
        RECT 131.420 55.380 134.930 55.430 ;
        RECT 140.100 55.380 141.060 56.980 ;
        RECT 147.120 55.400 148.080 55.460 ;
        RECT 142.600 55.380 148.080 55.400 ;
        RECT 131.420 54.470 148.080 55.380 ;
        RECT 133.400 54.440 148.080 54.470 ;
        RECT 133.400 54.420 144.300 54.440 ;
        RECT 130.105 45.230 130.435 46.285 ;
        RECT 132.760 45.230 133.080 53.530 ;
        RECT 133.400 45.230 134.360 54.420 ;
        RECT 137.180 54.400 138.260 54.420 ;
        RECT 141.330 54.400 142.410 54.420 ;
        RECT 143.340 53.570 144.300 54.420 ;
        RECT 147.120 54.380 148.080 54.440 ;
        RECT 135.320 51.260 136.280 53.530 ;
        RECT 130.055 44.900 133.080 45.230 ;
        RECT 108.720 42.620 127.370 43.820 ;
        RECT 108.630 32.400 109.950 33.600 ;
        RECT 126.170 32.410 127.370 42.620 ;
        RECT 132.750 41.630 133.080 44.900 ;
        RECT 133.390 41.630 134.360 45.230 ;
        RECT 132.760 41.120 133.080 41.630 ;
        RECT 133.400 41.120 134.360 41.630 ;
        RECT 132.750 40.520 133.080 41.120 ;
        RECT 132.750 37.520 133.070 40.520 ;
        RECT 133.390 39.250 134.360 41.120 ;
        RECT 135.310 49.930 136.280 51.260 ;
        RECT 135.310 49.420 136.270 49.930 ;
        RECT 135.310 45.820 136.280 49.420 ;
        RECT 133.390 37.520 134.350 39.250 ;
        RECT 135.310 35.340 136.270 45.820 ;
        RECT 139.975 45.270 140.305 45.300 ;
        RECT 142.670 45.270 142.990 53.570 ;
        RECT 143.310 52.230 144.300 53.570 ;
        RECT 143.310 51.030 144.270 52.230 ;
        RECT 139.965 44.940 142.990 45.270 ;
        RECT 139.975 44.910 140.305 44.940 ;
        RECT 142.660 41.670 142.990 44.940 ;
        RECT 142.670 41.160 142.990 41.670 ;
        RECT 142.660 40.690 142.990 41.160 ;
        RECT 143.300 49.970 144.270 51.030 ;
        RECT 143.300 49.460 144.260 49.970 ;
        RECT 143.300 45.860 144.270 49.460 ;
        RECT 142.660 37.560 142.980 40.690 ;
        RECT 143.300 37.560 144.260 45.860 ;
        RECT 145.230 45.270 146.190 53.570 ;
        RECT 145.220 41.670 146.190 45.270 ;
        RECT 145.230 41.160 146.190 41.670 ;
        RECT 145.220 39.630 146.190 41.160 ;
        RECT 145.220 35.690 146.180 39.630 ;
        RECT 150.810 38.000 151.770 95.250 ;
        RECT 150.810 35.690 151.900 38.000 ;
        RECT 132.760 35.290 136.350 35.340 ;
        RECT 132.760 35.020 143.000 35.290 ;
        RECT 97.630 23.120 98.590 26.720 ;
        RECT 98.910 23.120 99.870 29.360 ;
        RECT 97.750 21.310 98.590 23.120 ;
        RECT 103.150 20.720 104.470 22.780 ;
        RECT 85.935 19.170 92.990 20.370 ;
        RECT 103.090 19.400 104.530 20.720 ;
        RECT 85.935 17.605 88.985 19.170 ;
        RECT 17.920 13.460 19.920 13.490 ;
        RECT 17.920 11.460 24.850 13.460 ;
        RECT 71.240 12.555 72.440 17.605 ;
        RECT 69.995 11.800 73.045 12.555 ;
        RECT 77.965 11.800 81.015 12.555 ;
        RECT 85.935 11.800 88.985 12.555 ;
        RECT 91.790 11.800 92.990 19.170 ;
        RECT 108.690 16.630 109.890 32.400 ;
        RECT 132.760 29.760 133.080 35.020 ;
        RECT 135.310 34.970 143.000 35.020 ;
        RECT 135.310 33.360 136.270 34.970 ;
        RECT 133.400 27.660 134.360 33.360 ;
        RECT 135.310 31.360 136.280 33.360 ;
        RECT 135.320 29.760 136.280 31.360 ;
        RECT 142.680 29.750 143.000 34.970 ;
        RECT 145.220 34.730 159.400 35.690 ;
        RECT 145.220 33.350 146.180 34.730 ;
        RECT 143.320 27.780 144.280 33.350 ;
        RECT 145.220 31.480 146.200 33.350 ;
        RECT 145.240 29.750 146.200 31.480 ;
        RECT 106.980 16.080 107.540 16.140 ;
        RECT 108.690 16.080 132.550 16.630 ;
        RECT 106.980 15.520 132.550 16.080 ;
        RECT 106.980 15.460 107.540 15.520 ;
        RECT 108.690 15.430 132.550 15.520 ;
        RECT 17.920 11.430 19.920 11.460 ;
        RECT 69.995 10.600 92.990 11.800 ;
        RECT 69.995 9.505 73.045 10.600 ;
        RECT 77.965 9.505 81.015 10.600 ;
        RECT 85.935 9.505 88.985 10.600 ;
      LAYER met2 ;
        RECT 21.050 223.220 27.875 223.520 ;
        RECT 19.540 220.950 144.130 220.960 ;
        RECT 19.540 220.670 144.165 220.950 ;
        RECT 19.540 220.660 144.130 220.670 ;
        RECT 94.160 220.100 94.440 220.135 ;
        RECT 20.360 219.800 94.450 220.100 ;
        RECT 94.160 219.765 94.440 219.800 ;
        RECT 91.400 219.380 91.680 219.415 ;
        RECT 14.210 219.080 91.690 219.380 ;
        RECT 91.400 219.045 91.680 219.080 ;
        RECT 15.880 218.760 16.180 218.790 ;
        RECT 15.880 218.460 138.595 218.760 ;
        RECT 15.880 218.430 16.180 218.460 ;
        RECT 12.860 217.780 88.930 217.790 ;
        RECT 12.860 217.500 88.965 217.780 ;
        RECT 12.860 217.490 88.930 217.500 ;
        RECT 3.485 213.080 58.600 213.100 ;
        RECT 3.460 211.295 58.600 213.080 ;
        RECT 3.460 211.080 6.360 211.295 ;
        RECT 3.485 211.060 5.435 211.080 ;
        RECT 100.780 204.270 101.740 204.300 ;
        RECT 100.780 203.310 105.625 204.270 ;
        RECT 100.780 203.280 101.740 203.310 ;
        RECT 94.975 195.810 101.770 196.770 ;
        RECT 94.900 188.690 102.100 189.890 ;
        RECT 105.100 189.500 149.600 190.190 ;
        RECT 105.100 188.990 149.610 189.500 ;
        RECT 80.220 186.450 80.540 188.495 ;
        RECT 94.900 186.450 96.100 188.690 ;
        RECT 80.190 186.130 80.570 186.450 ;
        RECT 89.190 186.130 96.100 186.450 ;
        RECT 22.660 169.730 50.590 170.030 ;
        RECT 20.360 168.280 22.150 168.580 ;
        RECT 20.590 165.680 21.470 166.020 ;
        RECT 23.290 165.680 24.170 166.020 ;
        RECT 94.900 164.690 96.100 186.130 ;
        RECT 105.100 186.450 106.300 188.990 ;
        RECT 120.460 186.450 120.780 188.495 ;
        RECT 105.100 186.130 111.810 186.450 ;
        RECT 120.430 186.130 120.810 186.450 ;
        RECT 105.100 185.790 106.300 186.130 ;
        RECT 148.400 176.100 149.610 188.990 ;
        RECT 148.400 175.090 159.130 176.100 ;
        RECT 148.590 175.080 159.130 175.090 ;
        RECT 97.340 166.450 97.660 166.480 ;
        RECT 97.340 166.130 98.705 166.450 ;
        RECT 97.340 166.100 97.660 166.130 ;
        RECT 77.650 164.390 104.650 164.690 ;
        RECT 20.590 163.280 21.470 163.620 ;
        RECT 23.290 163.280 24.170 163.620 ;
        RECT 26.270 162.680 49.600 163.000 ;
        RECT 20.590 160.880 21.470 161.220 ;
        RECT 23.290 160.880 24.170 161.220 ;
        RECT 18.430 160.700 18.730 160.730 ;
        RECT 14.220 160.400 18.730 160.700 ;
        RECT 18.430 160.370 18.730 160.400 ;
        RECT 77.400 160.150 78.600 160.180 ;
        RECT 20.590 159.280 21.470 159.620 ;
        RECT 23.290 159.280 24.170 159.620 ;
        RECT 77.400 158.950 85.445 160.150 ;
        RECT 77.400 158.920 78.600 158.950 ;
        RECT 94.160 158.340 94.440 158.375 ;
        RECT 92.620 158.040 94.450 158.340 ;
        RECT 20.590 157.680 21.470 158.020 ;
        RECT 94.160 158.005 94.440 158.040 ;
        RECT 26.145 157.530 26.480 157.560 ;
        RECT 32.690 157.530 33.650 157.870 ;
        RECT 19.220 157.180 19.520 157.210 ;
        RECT 12.880 156.880 19.520 157.180 ;
        RECT 26.145 157.195 33.650 157.530 ;
        RECT 26.145 157.165 26.480 157.195 ;
        RECT 19.220 156.850 19.520 156.880 ;
        RECT 32.690 156.850 33.650 157.195 ;
        RECT 20.590 156.080 21.470 156.420 ;
        RECT 23.290 156.080 24.170 156.420 ;
        RECT 20.590 154.480 21.470 154.820 ;
        RECT 23.290 154.480 24.170 154.820 ;
        RECT 26.030 154.390 26.330 154.420 ;
        RECT 26.030 154.090 29.850 154.390 ;
        RECT 26.030 154.060 26.330 154.090 ;
        RECT 20.590 152.880 21.470 153.220 ;
        RECT 23.290 152.880 24.170 153.220 ;
        RECT 18.310 152.780 18.610 152.810 ;
        RECT 15.850 152.480 18.610 152.780 ;
        RECT 18.310 152.450 18.610 152.480 ;
        RECT 20.590 151.280 21.470 151.620 ;
        RECT 23.290 151.280 24.170 151.620 ;
        RECT 94.900 150.890 96.100 164.390 ;
        RECT 106.320 159.570 107.280 159.600 ;
        RECT 106.320 158.610 109.125 159.570 ;
        RECT 106.320 158.580 107.280 158.610 ;
        RECT 108.220 157.340 109.100 157.680 ;
        RECT 110.920 157.340 111.800 157.680 ;
        RECT 107.390 155.940 107.750 156.240 ;
        RECT 110.920 156.205 113.470 156.230 ;
        RECT 107.420 154.440 107.720 155.940 ;
        RECT 110.900 155.375 113.470 156.205 ;
        RECT 110.920 155.350 113.470 155.375 ;
        RECT 107.420 154.140 113.650 154.440 ;
        RECT 106.850 153.940 107.150 153.970 ;
        RECT 102.850 153.830 107.150 153.940 ;
        RECT 20.590 150.480 21.470 150.820 ;
        RECT 23.290 150.480 24.170 150.820 ;
        RECT 90.370 149.690 96.100 150.890 ;
        RECT 102.720 153.640 107.150 153.830 ;
        RECT 20.590 141.555 21.470 141.580 ;
        RECT 20.570 140.725 21.490 141.555 ;
        RECT 4.025 139.980 5.975 140.000 ;
        RECT 4.000 137.980 8.190 139.980 ;
        RECT 20.590 138.500 21.470 140.725 ;
        RECT 4.025 137.960 5.975 137.980 ;
        RECT 102.720 136.300 103.040 153.640 ;
        RECT 106.850 153.610 107.150 153.640 ;
        RECT 107.400 152.240 108.280 152.580 ;
        RECT 110.100 152.240 110.980 152.580 ;
        RECT 105.600 151.340 106.480 151.380 ;
        RECT 105.600 151.040 107.100 151.340 ;
        RECT 106.800 148.140 107.100 151.040 ;
        RECT 110.100 149.840 110.980 150.180 ;
        RECT 107.400 149.040 108.280 149.380 ;
        RECT 111.900 148.140 112.780 148.180 ;
        RECT 106.800 147.840 112.780 148.140 ;
        RECT 107.400 146.640 108.280 146.980 ;
        RECT 110.100 146.640 110.980 146.980 ;
        RECT 107.400 145.040 108.280 145.380 ;
        RECT 110.100 145.040 110.980 145.380 ;
        RECT 107.400 142.640 108.280 142.980 ;
        RECT 110.100 142.640 110.980 142.980 ;
        RECT 107.400 140.240 108.280 140.580 ;
        RECT 110.100 140.240 110.980 140.580 ;
        RECT 113.350 139.940 113.650 154.140 ;
        RECT 142.400 152.390 143.600 152.420 ;
        RECT 140.355 151.190 143.600 152.390 ;
        RECT 142.400 151.160 143.600 151.190 ;
        RECT 112.320 139.640 113.650 139.940 ;
        RECT 107.400 138.640 108.280 138.980 ;
        RECT 110.100 138.640 110.980 138.980 ;
        RECT 110.100 137.840 110.980 138.180 ;
        RECT 49.220 135.980 103.040 136.300 ;
        RECT 107.400 136.240 108.280 136.580 ;
        RECT 110.100 136.240 110.980 136.580 ;
        RECT 50.260 135.560 50.560 135.590 ;
        RECT 50.260 135.260 101.130 135.560 ;
        RECT 50.260 135.230 50.560 135.260 ;
        RECT 100.830 132.040 101.130 135.260 ;
        RECT 102.720 133.090 103.040 135.980 ;
        RECT 105.760 135.400 106.120 135.700 ;
        RECT 107.400 135.440 108.280 135.780 ;
        RECT 110.100 135.440 110.980 135.780 ;
        RECT 102.650 132.640 103.100 133.090 ;
        RECT 105.790 132.040 106.090 135.400 ;
        RECT 107.400 134.640 108.280 134.980 ;
        RECT 110.100 134.640 110.980 134.980 ;
        RECT 107.920 133.030 108.880 133.060 ;
        RECT 107.920 132.070 111.825 133.030 ;
        RECT 107.920 132.040 108.880 132.070 ;
        RECT 100.830 131.740 106.090 132.040 ;
        RECT 108.210 131.715 109.090 131.740 ;
        RECT 108.190 130.885 109.110 131.715 ;
        RECT 108.210 129.010 109.090 130.885 ;
        RECT 32.660 111.920 159.450 112.880 ;
        RECT 28.750 110.945 86.245 110.970 ;
        RECT 28.750 109.775 86.265 110.945 ;
        RECT 28.750 109.750 86.245 109.775 ;
        RECT 4.555 103.800 6.505 103.820 ;
        RECT 4.530 101.800 33.000 103.800 ;
        RECT 4.555 101.780 6.505 101.800 ;
        RECT 104.205 55.965 104.595 56.295 ;
        RECT 88.120 54.100 89.340 54.130 ;
        RECT 58.760 54.010 59.080 54.015 ;
        RECT 55.910 53.690 59.080 54.010 ;
        RECT 58.760 53.645 59.080 53.690 ;
        RECT 85.005 52.880 89.340 54.100 ;
        RECT 88.120 52.850 89.340 52.880 ;
        RECT 27.755 51.935 63.370 52.265 ;
        RECT 27.755 48.770 28.085 51.935 ;
        RECT 37.785 50.995 58.765 51.325 ;
        RECT 37.785 49.455 38.115 50.995 ;
        RECT 27.725 48.440 28.115 48.770 ;
        RECT 52.550 43.580 53.570 44.540 ;
        RECT 52.580 41.925 53.540 43.580 ;
        RECT 58.435 34.565 58.765 50.995 ;
        RECT 63.040 48.865 63.370 51.935 ;
        RECT 104.235 46.255 104.565 55.965 ;
        RECT 111.115 50.485 111.445 82.105 ;
        RECT 111.115 50.155 140.305 50.485 ;
        RECT 102.070 45.925 130.465 46.255 ;
        RECT 139.975 45.270 140.305 50.155 ;
        RECT 139.945 44.940 140.335 45.270 ;
        RECT 58.435 34.235 64.875 34.565 ;
        RECT 60.035 33.370 61.950 33.690 ;
        RECT 98.910 29.330 99.870 31.415 ;
        RECT 98.880 28.370 99.900 29.330 ;
        RECT 103.150 22.750 104.470 24.735 ;
        RECT 103.120 21.430 104.500 22.750 ;
        RECT 12.855 13.460 14.805 13.480 ;
        RECT 12.830 11.460 19.950 13.460 ;
        RECT 12.855 11.440 14.805 11.460 ;
      LAYER met3 ;
        RECT 143.790 224.200 144.170 224.520 ;
        RECT 88.590 223.710 88.970 224.030 ;
        RECT 27.525 223.520 27.855 223.545 ;
        RECT 31.060 223.520 31.440 223.530 ;
        RECT 27.525 223.220 31.440 223.520 ;
        RECT 27.525 223.195 27.855 223.220 ;
        RECT 31.060 223.210 31.440 223.220 ;
        RECT 88.630 217.805 88.930 223.710 ;
        RECT 91.350 223.640 91.730 223.960 ;
        RECT 94.110 223.720 94.490 224.040 ;
        RECT 91.390 219.395 91.690 223.640 ;
        RECT 94.150 220.115 94.450 223.720 ;
        RECT 138.250 223.650 138.570 224.030 ;
        RECT 94.135 219.785 94.465 220.115 ;
        RECT 91.375 219.065 91.705 219.395 ;
        RECT 138.260 218.785 138.560 223.650 ;
        RECT 143.830 220.975 144.130 224.200 ;
        RECT 143.815 220.645 144.145 220.975 ;
        RECT 138.245 218.435 138.575 218.785 ;
        RECT 88.615 217.475 88.945 217.805 ;
        RECT 0.980 213.080 3.040 213.130 ;
        RECT 0.980 211.080 5.460 213.080 ;
        RECT 0.980 211.020 3.040 211.080 ;
        RECT 3.940 141.380 6.370 143.710 ;
        RECT 4.000 137.980 6.000 141.380 ;
        RECT 20.590 140.700 21.470 167.030 ;
        RECT 23.290 150.230 24.170 213.100 ;
        RECT 80.195 188.470 80.565 188.475 ;
        RECT 94.900 188.470 96.100 196.890 ;
        RECT 80.195 188.150 96.100 188.470 ;
        RECT 80.195 188.145 80.565 188.150 ;
        RECT 84.225 160.150 85.425 160.175 ;
        RECT 94.900 160.150 96.100 188.150 ;
        RECT 104.645 188.870 105.605 204.295 ;
        RECT 104.645 187.910 124.180 188.870 ;
        RECT 98.355 166.450 98.685 166.475 ;
        RECT 98.340 166.130 101.160 166.450 ;
        RECT 98.355 166.105 98.685 166.130 ;
        RECT 100.840 164.690 101.160 166.130 ;
        RECT 84.225 158.950 96.100 160.150 ;
        RECT 97.600 159.290 103.000 164.690 ;
        RECT 84.225 158.925 85.425 158.950 ;
        RECT 94.135 158.340 94.465 158.355 ;
        RECT 96.440 158.340 96.760 158.380 ;
        RECT 94.135 158.040 96.760 158.340 ;
        RECT 94.135 158.025 94.465 158.040 ;
        RECT 96.440 158.000 96.760 158.040 ;
        RECT 108.145 155.170 109.105 159.595 ;
        RECT 110.920 155.350 111.800 158.690 ;
        RECT 108.145 154.730 110.680 155.170 ;
        RECT 108.145 154.210 110.980 154.730 ;
        RECT 107.400 131.740 108.280 153.590 ;
        RECT 110.100 134.390 110.980 154.210 ;
        RECT 123.220 151.490 124.180 187.910 ;
        RECT 140.375 152.390 141.575 152.415 ;
        RECT 120.500 146.090 125.900 151.490 ;
        RECT 128.300 146.090 133.700 151.490 ;
        RECT 138.370 151.190 141.575 152.390 ;
        RECT 140.375 151.165 141.575 151.190 ;
        RECT 123.000 143.690 123.400 146.090 ;
        RECT 130.800 143.690 131.200 146.090 ;
        RECT 120.500 140.270 125.900 143.690 ;
        RECT 116.020 139.310 125.900 140.270 ;
        RECT 110.845 133.030 111.805 133.055 ;
        RECT 116.020 133.030 116.980 139.310 ;
        RECT 120.500 138.790 125.900 139.310 ;
        RECT 128.300 138.790 133.700 143.690 ;
        RECT 120.500 138.290 133.700 138.790 ;
        RECT 110.845 132.070 116.980 133.030 ;
        RECT 110.845 132.045 111.805 132.070 ;
        RECT 107.400 130.860 109.090 131.740 ;
        RECT 0.930 103.800 3.360 103.980 ;
        RECT 0.930 101.800 6.530 103.800 ;
        RECT 0.930 101.650 3.360 101.800 ;
        RECT 58.735 53.665 59.105 53.995 ;
        RECT 52.555 41.945 53.565 42.905 ;
        RECT 52.580 37.490 53.540 41.945 ;
        RECT 50.670 32.090 56.070 37.490 ;
        RECT 58.760 33.690 59.080 53.665 ;
        RECT 85.025 52.855 86.245 110.970 ;
        RECT 102.090 46.255 102.420 46.280 ;
        RECT 100.595 45.900 102.420 46.255 ;
        RECT 100.595 43.080 100.925 45.900 ;
        RECT 98.190 37.680 103.590 43.080 ;
        RECT 60.055 33.690 60.385 33.715 ;
        RECT 58.380 33.370 60.385 33.690 ;
        RECT 58.760 33.340 59.080 33.370 ;
        RECT 60.055 33.345 60.385 33.370 ;
        RECT 98.910 31.395 99.870 37.680 ;
        RECT 98.885 30.435 99.895 31.395 ;
        RECT 103.150 24.715 104.470 27.020 ;
        RECT 103.125 23.395 104.495 24.715 ;
        RECT 3.740 13.460 6.170 13.710 ;
        RECT 3.740 11.460 14.830 13.460 ;
        RECT 3.740 11.380 6.170 11.460 ;
      LAYER met4 ;
        RECT 138.610 224.850 138.740 225.180 ;
        RECT 138.110 224.760 138.310 224.850 ;
        RECT 138.610 224.760 138.850 224.850 ;
        RECT 30.670 224.340 30.970 224.760 ;
        RECT 33.430 224.370 33.730 224.760 ;
        RECT 36.190 224.380 36.490 224.760 ;
        RECT 38.950 224.390 39.250 224.760 ;
        RECT 41.710 224.380 42.010 224.760 ;
        RECT 44.470 224.350 44.770 224.760 ;
        RECT 47.230 224.420 47.530 224.760 ;
        RECT 49.990 224.570 50.290 224.760 ;
        RECT 49.990 224.355 50.300 224.570 ;
        RECT 30.670 223.900 30.970 224.040 ;
        RECT 33.430 223.900 33.730 224.070 ;
        RECT 36.190 223.900 36.490 224.080 ;
        RECT 38.950 223.900 39.250 224.090 ;
        RECT 41.710 223.900 42.010 224.080 ;
        RECT 44.470 223.900 44.770 224.050 ;
        RECT 47.230 223.900 47.530 224.120 ;
        RECT 49.990 223.900 50.300 224.045 ;
        RECT 88.630 224.035 88.930 224.760 ;
        RECT 30.670 223.600 50.300 223.900 ;
        RECT 88.615 223.705 88.945 224.035 ;
        RECT 91.390 223.965 91.690 224.760 ;
        RECT 94.150 224.045 94.450 224.760 ;
        RECT 91.375 223.635 91.705 223.965 ;
        RECT 94.135 223.715 94.465 224.045 ;
        RECT 138.110 223.630 138.850 224.760 ;
        RECT 143.830 224.525 144.130 224.760 ;
        RECT 143.815 224.195 144.145 224.525 ;
        RECT 30.710 223.090 31.920 223.600 ;
        RECT 97.600 159.290 103.000 164.690 ;
        RECT 96.435 158.340 96.765 158.355 ;
        RECT 99.050 158.340 99.350 159.290 ;
        RECT 96.435 158.040 99.350 158.340 ;
        RECT 96.435 158.025 96.765 158.040 ;
        RECT 120.500 146.090 125.900 151.490 ;
        RECT 128.300 150.390 133.700 151.490 ;
        RECT 138.395 150.390 139.595 152.395 ;
        RECT 128.300 149.190 139.595 150.390 ;
        RECT 128.300 146.090 133.700 149.190 ;
        RECT 123.000 143.690 123.400 146.090 ;
        RECT 130.800 143.690 131.200 146.090 ;
        RECT 120.500 138.790 125.900 143.690 ;
        RECT 128.300 138.790 133.700 143.690 ;
        RECT 120.500 138.290 133.700 138.790 ;
        RECT 98.190 37.680 103.590 43.080 ;
        RECT 102.210 37.620 103.260 37.680 ;
        RECT 102.265 37.550 103.220 37.620 ;
        RECT 50.670 33.690 56.070 37.490 ;
        RECT 58.405 33.690 58.735 33.695 ;
        RECT 50.670 33.370 58.735 33.690 ;
        RECT 50.670 32.090 56.070 33.370 ;
        RECT 58.405 33.365 58.735 33.370 ;
        RECT 102.265 31.215 103.215 37.550 ;
        RECT 102.265 30.265 104.085 31.215 ;
        RECT 103.135 27.290 104.085 30.265 ;
        RECT 103.135 26.980 104.520 27.290 ;
        RECT 103.135 25.675 104.475 26.980 ;
        RECT 103.135 25.625 104.085 25.675 ;
  END
END tt_um_jnw_wulffern
END LIBRARY

